-------------------------------------------------------------------------------
-- Title      : Cpix detector conversion look-up table package
-------------------------------------------------------------------------------
-- File       : CpixLUT.vhd
-- Author     : Maciej Kwiatkowski <mkwiatko@slac.stanford.edu>
-- Company    : SLAC National Accelerator Laboratory
-- Created    : 03/09/2016
-- Last update: 03/09/2016
-- Platform   : Vivado 2014.4
-- Standard   : VHDL'93/02
-------------------------------------------------------------------------------
-- Description: Cpix detector conversion look-up table package
-------------------------------------------------------------------------------
-- This file is part of 'CPIX Development Firmware'.
-- It is subject to the license terms in the LICENSE.txt file found in the 
-- top-level directory of this distribution and at: 
--    https://confluence.slac.stanford.edu/display/ppareg/LICENSE.html. 
-- No part of 'CPIX Development Firmware', including this file, 
-- may be copied, modified, propagated, or distributed except according to 
-- the terms contained in the LICENSE.txt file.
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package CpixLUTPkg is
   
   type NatArray is array (natural range <>) of natural;
   constant CPIX_NORMAL_SIM_ARRAY_C : NatArray(0 to 32767) := (
      0 ,1 ,240 ,2 ,15345 ,241 ,1023 ,3 ,20898 ,15346 ,7775 ,242 ,480 ,1024 ,3840 ,4 ,1263 ,20899 ,20038 ,15347 ,28380 ,7776 ,18061 ,243 ,9120 ,481 ,29558 ,1025 ,26919 ,3841 ,15585 ,5 ,31160 ,1264 ,5052 ,20900 ,16151 ,20039 ,720 ,15348 ,4080 ,28381 ,16368 ,7777 ,11065 ,18062 ,9546 ,244 ,30690 ,9121 ,21581 ,482 ,8015 ,29559 ,7432 ,1026 ,10194 ,26920 ,21138 ,3842 ,2046 ,15586 ,10455 ,6 ,16502 ,31161 ,19185 ,1265 ,29798 ,5053 ,12444 ,20901 ,8798 ,16152 ,9360 ,20040 ,30543 ,721 ,22195 ,15349 ,24564 ,4081 ,13956 ,28382 ,1905 ,16369 ,27159 ,7778 ,15825 ,11066 ,18755 ,18063 ,23436 ,9547 ,21921 ,245 ,18301 ,30691 ,5606 ,9122 ,4863 ,21582 ,24026 ,483 ,6777 ,8016 ,26386 ,29560 ,3476 ,7433 ,28620 ,1027 ,5224 ,10195 ,1503 ,26921 ,19462 ,21139 ,23120 ,3843 ,8191 ,2047 ,2533 ,15587 ,20278 ,10456 ,127 ,7 ,7672 ,16503 ,13459 ,31162 ,2431 ,19186 ,26522 ,1266 ,9497 ,29799 ,6143 ,5054 ,19084 ,12445 ,8255 ,20902 ,10865 ,8799 ,30930 ,16153 ,18893 ,9361 ,24738 ,20041 ,14749 ,30544 ,29403 ,722 ,21821 ,22196 ,17020 ,15350 ,21061 ,24565 ,2992 ,4082 ,21378 ,13957 ,12136 ,28383 ,20376 ,1906 ,10434 ,16370 ,14095 ,27160 ,31659 ,7779 ,11615 ,15826 ,18393 ,11067 ,14684 ,18756 ,2286 ,18064 ,10695 ,23437 ,17605 ,9548 ,24465 ,21922 ,24062 ,246 ,9029 ,18302 ,27942 ,30692 ,28220 ,5607 ,11305 ,9123 ,9786 ,4864 ,24953 ,21583 ,15550 ,24027 ,2616 ,484 ,4212 ,6778 ,14618 ,8017 ,16608 ,26387 ,26099 ,29561 ,6698 ,3477 ,4320 ,7434 ,27299 ,28621 ,29848 ,1028 ,10958 ,5225 ,31400 ,10196 ,13876 ,1504 ,28071 ,26922 ,29704 ,19463 ,13563 ,21140 ,5292 ,23121 ,10143 ,3844 ,960 ,8192 ,28673 ,2048 ,31290 ,2534 ,24642 ,15588 ,30581 ,20279 ,639 ,10457 ,7680 ,128 ,16391 ,8 ,
      20271 ,7673 ,16895 ,16504 ,10569 ,13460 ,3716 ,31163 ,28860 ,2432 ,22036 ,19187 ,16703 ,26523 ,12321 ,1267 ,27111 ,9498 ,12088 ,29800 ,26626 ,6144 ,28736 ,5055 ,23878 ,19085 ,7017 ,12446 ,25539 ,8256 ,5484 ,20903 ,11386 ,10866 ,18541 ,8800 ,32598 ,30931 ,24335 ,16154 ,17391 ,18894 ,31267 ,9362 ,5846 ,24739 ,23237 ,20042 ,24266 ,14750 ,25800 ,30545 ,15050 ,29404 ,9895 ,723 ,23764 ,21822 ,21737 ,22197 ,4566 ,17021 ,5103 ,15351 ,23360 ,21062 ,10789 ,24566 ,27737 ,2993 ,28784 ,4083 ,3156 ,21379 ,17174 ,13958 ,28033 ,12137 ,19702 ,28384 ,30018 ,20377 ,5464 ,1907 ,21901 ,10435 ,17000 ,16371 ,25685 ,14096 ,22777 ,27161 ,1743 ,31660 ,2651 ,7780 ,26232 ,11616 ,17689 ,15827 ,2773 ,18394 ,32183 ,11068 ,32067 ,14685 ,8431 ,18757 ,7102 ,2287 ,4159 ,18065 ,6075 ,10696 ,32220 ,23438 ,13268 ,17606 ,20518 ,9549 ,367 ,24466 ,4780 ,21923 ,16902 ,24063 ,1927 ,247 ,631 ,9030 ,26832 ,18303 ,18995 ,27943 ,3388 ,30693 ,32131 ,28221 ,16065 ,5608 ,11684 ,11306 ,11217 ,9124 ,31496 ,9787 ,2199 ,4865 ,29267 ,24954 ,23676 ,21584 ,22161 ,15551 ,10109 ,24028 ,12287 ,2617 ,2111 ,485 ,27399 ,4213 ,3069 ,6779 ,13738 ,14619 ,12960 ,8018 ,25399 ,16609 ,8169 ,26388 ,30404 ,26100 ,2145 ,29562 ,23291 ,6699 ,24804 ,3478 ,11478 ,4321 ,26674 ,7435 ,25836 ,27300 ,7348 ,28622 ,14196 ,29849 ,20397 ,1029 ,22604 ,10959 ,16742 ,5226 ,27813 ,31401 ,22862 ,10197 ,21222 ,13877 ,5989 ,1505 ,19425 ,28072 ,6192 ,26923 ,12684 ,29705 ,22710 ,19464 ,20767 ,13564 ,31713 ,21141 ,11773 ,5293 ,30845 ,23122 ,11723 ,10144 ,30038 ,3845 ,19123 ,961 ,24891 ,8193 ,5402 ,28674 ,30783 ,2049 ,22435 ,31291 ,30759 ,2535 ,8455 ,24643 ,18249 ,15589 ,23369 ,30582 ,13587 ,20280 ,9600 ,640 ,22613 ,10458 ,26410 ,7681 ,9038 ,129 ,16511 ,16392 ,519 ,9 ,
      2040 ,20272 ,24459 ,7674 ,4560 ,16896 ,14190 ,16505 ,14852 ,10570 ,6938 ,13461 ,3349 ,3717 ,8304 ,31164 ,26029 ,28861 ,25306 ,2433 ,22944 ,22037 ,27539 ,19188 ,30088 ,16704 ,5698 ,26524 ,8630 ,12322 ,22797 ,1268 ,26339 ,27112 ,19991 ,9499 ,29356 ,12089 ,31353 ,29801 ,16018 ,26627 ,13540 ,6145 ,4733 ,28737 ,16848 ,5056 ,1434 ,23879 ,4452 ,19086 ,20569 ,7018 ,6450 ,12447 ,19778 ,25540 ,4405 ,8257 ,14858 ,5485 ,4899 ,20904 ,5393 ,11387 ,9269 ,10867 ,30353 ,18542 ,17878 ,8801 ,8892 ,32599 ,19825 ,30932 ,28182 ,24336 ,6549 ,16155 ,11545 ,17392 ,4665 ,18895 ,13246 ,31268 ,25171 ,9363 ,15207 ,5847 ,2928 ,24740 ,23536 ,23238 ,28460 ,20043 ,14979 ,24267 ,22497 ,14751 ,23843 ,25801 ,15790 ,30546 ,2856 ,15051 ,12660 ,29405 ,18593 ,9896 ,2233 ,724 ,31092 ,23765 ,15472 ,21823 ,25193 ,21738 ,25587 ,22198 ,14786 ,4567 ,10026 ,17022 ,10576 ,5104 ,27181 ,15352 ,952 ,23361 ,15271 ,21063 ,4007 ,10790 ,5532 ,24567 ,10383 ,27738 ,9712 ,2994 ,22122 ,28785 ,31585 ,4084 ,29488 ,3157 ,12213 ,21380 ,13803 ,17175 ,8964 ,13959 ,15753 ,28034 ,29944 ,12138 ,13386 ,19703 ,9821 ,28385 ,18230 ,30019 ,11198 ,20378 ,23218 ,5465 ,19683 ,1908 ,28601 ,21902 ,3821 ,10436 ,31640 ,17001 ,2597 ,16372 ,28311 ,25686 ,31566 ,14097 ,16829 ,22778 ,6530 ,27162 ,18821 ,1744 ,14905 ,31661 ,6944 ,2652 ,14116 ,7781 ,24882 ,26233 ,4946 ,11617 ,13048 ,17690 ,17525 ,15828 ,12888 ,2774 ,6604 ,18395 ,21545 ,32184 ,31530 ,11069 ,20208 ,32068 ,1200 ,14686 ,12754 ,8432 ,1371 ,18758 ,22532 ,7103 ,29158 ,2288 ,28913 ,4160 ,25705 ,18066 ,14024 ,6076 ,17969 ,10697 ,879 ,32221 ,12850 ,23439 ,8359 ,13269 ,30821 ,17607 ,12777 ,20519 ,28330 ,9550 ,15279 ,368 ,20790 ,24467 ,28109 ,4781 ,7920 ,21924 ,16631 ,16903 ,26840 ,24064 ,13467 ,1928 ,20951 ,248 ,
      2526 ,632 ,4773 ,9031 ,10019 ,26833 ,24176 ,18304 ,15700 ,18996 ,21455 ,27944 ,7309 ,3389 ,14924 ,30694 ,19632 ,32132 ,11855 ,28222 ,22311 ,16066 ,6247 ,5609 ,13121 ,11685 ,25950 ,11307 ,18633 ,11218 ,12494 ,9125 ,12817 ,31497 ,6497 ,9788 ,17845 ,2200 ,27506 ,4866 ,19291 ,29268 ,10935 ,24955 ,24143 ,23677 ,23710 ,21585 ,23993 ,22162 ,7399 ,15552 ,11272 ,10110 ,24705 ,24029 ,24302 ,12288 ,20485 ,2618 ,3355 ,2112 ,31680 ,486 ,22426 ,27400 ,32492 ,4214 ,31847 ,3070 ,14335 ,6780 ,31899 ,13739 ,13674 ,14620 ,4282 ,12961 ,9214 ,8019 ,17321 ,25400 ,19757 ,16610 ,10674 ,8170 ,23743 ,26389 ,3556 ,30405 ,20616 ,26101 ,1621 ,2146 ,1763 ,29563 ,4489 ,23292 ,21301 ,6700 ,3272 ,24805 ,7065 ,3479 ,30160 ,11479 ,27789 ,4322 ,3232 ,26675 ,18840 ,7436 ,12376 ,25837 ,8517 ,27301 ,1150 ,7349 ,12038 ,28623 ,25421 ,14197 ,24183 ,29850 ,3723 ,20398 ,21618 ,1030 ,24634 ,22605 ,7912 ,10960 ,31963 ,16743 ,21480 ,5227 ,27685 ,27814 ,5886 ,31402 ,13699 ,22863 ,29301 ,10198 ,26762 ,21223 ,5911 ,13878 ,7142 ,5990 ,23926 ,1506 ,15014 ,19426 ,6347 ,28073 ,25049 ,6193 ,2671 ,26924 ,17250 ,12685 ,27019 ,29706 ,19850 ,22711 ,19324 ,19465 ,8495 ,20768 ,1481 ,13565 ,14295 ,31714 ,6963 ,21142 ,6629 ,11774 ,28986 ,5294 ,6383 ,30846 ,30444 ,23123 ,17342 ,11724 ,9737 ,10145 ,8310 ,30039 ,15651 ,3846 ,18240 ,19124 ,16090 ,962 ,29643 ,24892 ,14034 ,8194 ,6014 ,5403 ,14989 ,28675 ,26349 ,30784 ,14135 ,2050 ,5332 ,22436 ,4499 ,31292 ,12827 ,30760 ,22061 ,2536 ,17260 ,8456 ,22250 ,24644 ,17199 ,18250 ,24988 ,15590 ,24978 ,23370 ,26242 ,30583 ,11396 ,13588 ,1333 ,20281 ,27409 ,9601 ,6168 ,641 ,3516 ,22614 ,19133 ,10459 ,21071 ,26411 ,11105 ,7682 ,9385 ,9039 ,10968 ,130 ,3895 ,16512 ,18311 ,16393 ,31170 ,520 ,7800 ,10 ,
      26914 ,2041 ,23431 ,20273 ,21816 ,24460 ,27294 ,7675 ,25534 ,4561 ,1738 ,16897 ,12282 ,14191 ,11718 ,16506 ,8625 ,14853 ,23531 ,10571 ,13381 ,6939 ,28908 ,13462 ,18628 ,3350 ,1616 ,3718 ,25044 ,8305 ,17194 ,31165 ,25039 ,26030 ,25488 ,28862 ,7588 ,25307 ,13154 ,2434 ,10303 ,22945 ,26076 ,22038 ,25266 ,27540 ,13822 ,19189 ,29089 ,30089 ,32455 ,16705 ,25085 ,5699 ,14436 ,26525 ,20637 ,8631 ,30232 ,12323 ,26035 ,22798 ,7856 ,1269 ,19416 ,26340 ,8752 ,27113 ,434 ,19992 ,30644 ,9500 ,2385 ,29357 ,10649 ,12090 ,7634 ,31354 ,8983 ,29802 ,29221 ,16019 ,25353 ,26628 ,8409 ,13541 ,12638 ,6146 ,2727 ,4734 ,25639 ,28738 ,25493 ,16849 ,11340 ,5057 ,6337 ,1435 ,27639 ,23880 ,26303 ,4453 ,21025 ,19087 ,31801 ,20570 ,25375 ,7019 ,3309 ,6451 ,2480 ,12448 ,13200 ,19779 ,2810 ,25541 ,4687 ,4406 ,25983 ,8258 ,23172 ,14859 ,15707 ,5486 ,28867 ,4900 ,13978 ,20905 ,13868 ,5394 ,871 ,11388 ,32682 ,9270 ,18666 ,10868 ,30493 ,30354 ,13649 ,18543 ,27072 ,17879 ,12232 ,8802 ,3628 ,8893 ,15118 ,32600 ,1819 ,19826 ,20701 ,30933 ,30316 ,28183 ,7220 ,24337 ,7593 ,6550 ,19235 ,16156 ,26752 ,11546 ,27586 ,17393 ,16284 ,4666 ,11924 ,18896 ,11457 ,13247 ,7994 ,31269 ,16808 ,25172 ,11251 ,9364 ,6875 ,15208 ,25887 ,5848 ,16305 ,2929 ,21674 ,24741 ,9931 ,23537 ,32371 ,23239 ,25312 ,28461 ,21399 ,20044 ,5980 ,14980 ,30126 ,24268 ,10349 ,22498 ,15984 ,14752 ,3122 ,23844 ,22401 ,25802 ,20864 ,15791 ,20342 ,30547 ,12550 ,2857 ,14552 ,15052 ,20185 ,12661 ,12527 ,29406 ,2351 ,18594 ,22991 ,9897 ,13159 ,2234 ,3176 ,725 ,23916 ,31093 ,28524 ,23766 ,32690 ,15473 ,22084 ,21824 ,23025 ,25194 ,3045 ,21739 ,1394 ,25588 ,29507 ,22199 ,4015 ,14787 ,31736 ,4568 ,8083 ,10027 ,31971 ,17023 ,26122 ,10577 ,19003 ,5105 ,2439 ,27182 ,9158 ,15353 ,
      5217 ,953 ,6068 ,23362 ,31085 ,15272 ,12369 ,21064 ,13193 ,4008 ,12013 ,10791 ,25761 ,5533 ,29963 ,24568 ,17124 ,10384 ,9662 ,27739 ,19557 ,9713 ,11963 ,2995 ,30278 ,22123 ,19916 ,28786 ,10308 ,31586 ,28255 ,4085 ,31953 ,29489 ,15966 ,3158 ,20683 ,12214 ,11906 ,21381 ,14418 ,13804 ,27276 ,17176 ,12620 ,8965 ,21007 ,13960 ,27470 ,15754 ,12924 ,28035 ,11945 ,29945 ,11888 ,12139 ,7513 ,13387 ,8677 ,19704 ,22950 ,9822 ,12157 ,28386 ,22595 ,18231 ,22844 ,30020 ,23658 ,11199 ,12942 ,20379 ,9877 ,23219 ,3698 ,5466 ,16982 ,19684 ,32165 ,1909 ,23102 ,28602 ,12426 ,21903 ,18043 ,3822 ,702 ,10437 ,2268 ,31641 ,26504 ,17002 ,26081 ,2598 ,28053 ,16373 ,7902 ,28312 ,17507 ,25687 ,8946 ,31567 ,19665 ,14098 ,6432 ,16830 ,14172 ,22779 ,25153 ,6531 ,15772 ,27163 ,12020 ,18822 ,14317 ,1745 ,6229 ,14906 ,27488 ,31662 ,30426 ,6945 ,21462 ,2653 ,22043 ,14117 ,1315 ,7782 ,31392 ,24883 ,17961 ,26234 ,28516 ,4947 ,8695 ,11618 ,18489 ,13049 ,21276 ,17691 ,5807 ,17526 ,26571 ,15829 ,14482 ,12889 ,14517 ,2775 ,30999 ,6605 ,6280 ,18396 ,30895 ,21546 ,22675 ,32185 ,25271 ,31531 ,19722 ,11070 ,27675 ,20209 ,19363 ,32069 ,1843 ,1201 ,27237 ,14687 ,3210 ,12755 ,3454 ,8433 ,25131 ,1372 ,13405 ,18759 ,31023 ,22533 ,5745 ,7104 ,13319 ,29159 ,7531 ,2289 ,3577 ,28914 ,19581 ,4161 ,27545 ,25706 ,5642 ,18067 ,22853 ,14025 ,22335 ,6077 ,24374 ,17970 ,22344 ,10698 ,7166 ,880 ,30135 ,32222 ,8761 ,12851 ,9840 ,23440 ,16235 ,8360 ,23609 ,13270 ,29135 ,30822 ,22968 ,17608 ,17796 ,12778 ,12999 ,20520 ,13827 ,28331 ,10520 ,9551 ,29291 ,15280 ,4955 ,369 ,9278 ,20791 ,12175 ,24468 ,32501 ,28110 ,26650 ,4782 ,8852 ,7921 ,16099 ,21925 ,10798 ,16632 ,20107 ,16904 ,18917 ,26841 ,16751 ,24065 ,759 ,13468 ,27951 ,1929 ,19194 ,20952 ,28404 ,249 ,
      21132 ,2527 ,17599 ,633 ,21731 ,4774 ,7342 ,9032 ,4399 ,10020 ,14899 ,26834 ,20479 ,24177 ,9731 ,18305 ,30226 ,15701 ,32365 ,18997 ,8671 ,21456 ,19575 ,27945 ,32333 ,7310 ,32307 ,3390 ,29094 ,14925 ,575 ,30695 ,14285 ,19633 ,26472 ,32133 ,15934 ,11856 ,11981 ,28223 ,23577 ,22312 ,27919 ,16067 ,17929 ,6248 ,3422 ,5610 ,32423 ,13122 ,1584 ,11686 ,27607 ,25951 ,10617 ,11308 ,15086 ,18634 ,32339 ,11219 ,30094 ,12495 ,3013 ,9126 ,20758 ,12818 ,29126 ,31498 ,11166 ,6498 ,9680 ,9789 ,4633 ,17846 ,9994 ,2201 ,24427 ,27507 ,13508 ,4867 ,28954 ,19292 ,6315 ,29269 ,26210 ,10936 ,14957 ,24956 ,11823 ,24144 ,20453 ,23678 ,32460 ,23711 ,27757 ,21586 ,1471 ,23994 ,18723 ,22163 ,5020 ,7400 ,7743 ,15553 ,14586 ,11273 ,607 ,10111 ,13427 ,24706 ,10402 ,24030 ,25768 ,24303 ,6985 ,12289 ,17657 ,20486 ,17142 ,2619 ,2167 ,3356 ,7316 ,2113 ,16710 ,31681 ,30727 ,487 ,29696 ,22427 ,8351 ,27401 ,23017 ,32493 ,19934 ,4215 ,9446 ,31848 ,25925 ,3071 ,32028 ,14336 ,19029 ,6781 ,7246 ,31900 ,8567 ,13740 ,5783 ,13675 ,1983 ,14621 ,2891 ,4283 ,32397 ,12962 ,25090 ,9215 ,28804 ,8020 ,17240 ,17322 ,13101 ,25401 ,15187 ,19758 ,15733 ,16611 ,6678 ,10675 ,9100 ,8171 ,25665 ,23744 ,22141 ,26390 ,17776 ,3557 ,30258 ,30406 ,2707 ,20617 ,30296 ,26102 ,1642 ,1622 ,32313 ,2147 ,5704 ,1764 ,31211 ,29564 ,22701 ,4490 ,23600 ,23293 ,27866 ,21302 ,3764 ,6701 ,12584 ,3273 ,19607 ,24806 ,11029 ,7066 ,31604 ,3480 ,29024 ,30161 ,5159 ,11480 ,13025 ,27790 ,10326 ,4323 ,1662 ,3233 ,15908 ,26676 ,14441 ,18841 ,27977 ,7437 ,19314 ,12377 ,8703 ,25838 ,18674 ,8518 ,28273 ,27302 ,19942 ,1151 ,16041 ,7350 ,24842 ,12039 ,191 ,28624 ,5540 ,25422 ,18431 ,14198 ,17414 ,24184 ,21488 ,29851 ,18129 ,3724 ,3396 ,20399 ,26530 ,21619 ,4103 ,1031 ,
      23113 ,24635 ,20511 ,22606 ,25580 ,7913 ,12031 ,10961 ,25976 ,31964 ,27481 ,16744 ,17135 ,21481 ,16447 ,5228 ,3956 ,27686 ,31034 ,27815 ,14493 ,5887 ,24209 ,31403 ,16246 ,13700 ,4607 ,22864 ,20642 ,29302 ,10809 ,10199 ,6373 ,26763 ,6886 ,21224 ,3639 ,5912 ,16943 ,13879 ,12561 ,7143 ,9763 ,5991 ,29904 ,23927 ,4026 ,1507 ,29232 ,15015 ,16573 ,19427 ,22276 ,6348 ,13211 ,28074 ,1784 ,25050 ,29100 ,6194 ,8636 ,2672 ,18337 ,26925 ,11764 ,17251 ,17787 ,12686 ,7257 ,27020 ,10052 ,29707 ,29035 ,19851 ,24118 ,22712 ,2954 ,19325 ,5551 ,19466 ,28965 ,8496 ,4431 ,20769 ,18372 ,1482 ,25779 ,13566 ,5724 ,14296 ,32434 ,31715 ,30237 ,6964 ,16552 ,21143 ,28976 ,6630 ,14237 ,11775 ,29184 ,28987 ,29981 ,5295 ,17076 ,6384 ,29243 ,30847 ,3967 ,30445 ,26866 ,23124 ,29970 ,17343 ,27351 ,11725 ,11567 ,9738 ,16454 ,10146 ,29440 ,8311 ,14931 ,30040 ,12328 ,15652 ,24586 ,3847 ,10135 ,18241 ,28322 ,19125 ,29499 ,16091 ,183 ,963 ,20219 ,29644 ,7374 ,24893 ,21862 ,14035 ,15290 ,8195 ,11556 ,6015 ,24506 ,5404 ,30871 ,14990 ,31103 ,28676 ,31231 ,26350 ,1445 ,30785 ,26040 ,14136 ,9064 ,2051 ,17332 ,5333 ,21763 ,22437 ,21977 ,4500 ,12387 ,31293 ,7043 ,12828 ,24004 ,30761 ,19643 ,22062 ,7721 ,2537 ,27340 ,17261 ,6640 ,8457 ,26773 ,22251 ,4806 ,24645 ,5343 ,17200 ,581 ,18251 ,22803 ,24989 ,21082 ,15591 ,30029 ,24979 ,10511 ,23371 ,4346 ,26243 ,6086 ,30584 ,23477 ,11397 ,24277 ,13589 ,27122 ,1334 ,665 ,20282 ,29429 ,27410 ,23302 ,9602 ,31507 ,6169 ,20319 ,642 ,12695 ,3517 ,17631 ,22615 ,7861 ,19134 ,23380 ,10460 ,15641 ,21072 ,11626 ,26412 ,10876 ,11106 ,2559 ,7683 ,4223 ,9386 ,2087 ,9040 ,18781 ,10969 ,971 ,131 ,24575 ,3896 ,21164 ,16513 ,26960 ,18312 ,5235 ,16394 ,29584 ,31171 ,30701 ,521 ,1274 ,7801 ,71 ,11 ,
      476 ,26915 ,11061 ,2042 ,30539 ,23432 ,3472 ,20274 ,19080 ,21817 ,14091 ,24461 ,15546 ,27295 ,5288 ,7676 ,16699 ,25535 ,5842 ,4562 ,28029 ,1739 ,7098 ,16898 ,11680 ,12283 ,30400 ,14192 ,19421 ,11719 ,8451 ,16507 ,3345 ,8626 ,4729 ,14854 ,28178 ,23532 ,18589 ,10572 ,22118 ,13382 ,31636 ,6940 ,21541 ,28909 ,12773 ,13463 ,7305 ,18629 ,24139 ,3351 ,4278 ,1617 ,3228 ,3719 ,13695 ,25045 ,14291 ,8306 ,26345 ,17195 ,3512 ,31166 ,12278 ,25040 ,25262 ,26031 ,7630 ,25489 ,3305 ,28863 ,27068 ,7589 ,16804 ,25308 ,20860 ,13155 ,1390 ,2435 ,25757 ,10304 ,12616 ,22946 ,16978 ,26077 ,25149 ,22039 ,5803 ,25267 ,25127 ,27541 ,8757 ,13823 ,8848 ,19190 ,20475 ,29090 ,17925 ,30090 ,24423 ,32456 ,13423 ,16706 ,32024 ,25086 ,25661 ,5700 ,11025 ,14437 ,24838 ,26526 ,17131 ,20638 ,29900 ,8632 ,2950 ,30233 ,3963 ,12324 ,21858 ,26036 ,19639 ,22799 ,27118 ,7857 ,18777 ,1270 ,15542 ,19417 ,21537 ,26341 ,20856 ,8753 ,11021 ,27114 ,32724 ,435 ,3796 ,19993 ,32728 ,30645 ,1219 ,9501 ,5009 ,2386 ,9316 ,29358 ,18019 ,10650 ,1861 ,12091 ,2003 ,7635 ,23076 ,31355 ,439 ,8984 ,6733 ,29803 ,23983 ,29222 ,27898 ,16020 ,7973 ,25354 ,27255 ,26629 ,8148 ,8410 ,16347 ,13542 ,3800 ,12639 ,10914 ,6147 ,18712 ,2728 ,17561 ,4735 ,16326 ,25640 ,21334 ,28739 ,29755 ,25494 ,26478 ,16850 ,19997 ,11341 ,14705 ,5058 ,10100 ,6338 ,22666 ,1436 ,5182 ,27640 ,19381 ,23881 ,917 ,26304 ,18205 ,4454 ,32732 ,21026 ,23325 ,19088 ,14575 ,31802 ,8125 ,20571 ,28578 ,25376 ,11434 ,7020 ,15507 ,3310 ,23632 ,6452 ,30649 ,2481 ,32087 ,12449 ,24695 ,13201 ,18497 ,19780 ,30501 ,2811 ,4522 ,25542 ,9454 ,4688 ,5440 ,4407 ,1223 ,25984 ,20227 ,8259 ,10391 ,23173 ,22733 ,14860 ,13914 ,15708 ,27693 ,5487 ,14641 ,28868 ,32139 ,4901 ,9505 ,13979 ,323 ,20906 ,
      4856 ,13869 ,2766 ,5395 ,23836 ,872 ,3265 ,11389 ,26296 ,32683 ,8939 ,9271 ,5013 ,18667 ,29177 ,10869 ,24416 ,30494 ,1694 ,30355 ,3674 ,13650 ,13337 ,18544 ,8587 ,27073 ,14392 ,17880 ,2390 ,12233 ,10259 ,8803 ,17835 ,3629 ,827 ,8894 ,32556 ,15119 ,7549 ,32601 ,15164 ,1820 ,21355 ,19827 ,9320 ,20702 ,26708 ,30934 ,9983 ,30317 ,18959 ,28184 ,21695 ,7221 ,32646 ,24338 ,23800 ,7594 ,15940 ,6551 ,29362 ,19236 ,2307 ,16157 ,31487 ,26753 ,14473 ,11547 ,26190 ,27587 ,5763 ,17394 ,20165 ,16285 ,13361 ,4667 ,18023 ,11925 ,30979 ,18897 ,20747 ,11458 ,26606 ,13248 ,1885 ,7995 ,18873 ,31270 ,12734 ,16809 ,22924 ,25173 ,10654 ,11252 ,7122 ,9365 ,6487 ,6876 ,17463 ,15209 ,1701 ,25888 ,21999 ,5849 ,28558 ,16306 ,28009 ,2930 ,1865 ,21675 ,22551 ,24742 ,9669 ,9932 ,19872 ,23538 ,10747 ,32372 ,31041 ,23240 ,13760 ,25313 ,11862 ,28462 ,12095 ,21400 ,7469 ,20045 ,24945 ,5981 ,6596 ,14981 ,22393 ,30127 ,19599 ,24269 ,18197 ,10350 ,15246 ,22499 ,2007 ,15985 ,11512 ,14753 ,26199 ,3123 ,24233 ,23845 ,22571 ,22402 ,31463 ,25803 ,31127 ,20865 ,5191 ,15792 ,7639 ,20343 ,4179 ,30548 ,19281 ,12551 ,17743 ,2858 ,20725 ,14553 ,30193 ,15053 ,17299 ,20186 ,24542 ,12662 ,23080 ,12528 ,28932 ,29407 ,6304 ,2352 ,29056 ,18595 ,5947 ,22992 ,3595 ,9898 ,31920 ,13160 ,11987 ,2235 ,31359 ,3177 ,16202 ,726 ,23667 ,23917 ,6271 ,31094 ,31454 ,28525 ,24383 ,23767 ,23950 ,32691 ,10358 ,15474 ,443 ,22085 ,25724 ,21825 ,11812 ,23026 ,27875 ,25195 ,11175 ,3046 ,27563 ,21740 ,7266 ,1395 ,19531 ,25589 ,8988 ,29508 ,4355 ,22200 ,23700 ,4016 ,13057 ,14788 ,30362 ,31737 ,5660 ,4569 ,31856 ,8084 ,28760 ,10028 ,6737 ,31972 ,29652 ,17024 ,27746 ,26123 ,15864 ,10578 ,24762 ,19004 ,27822 ,5106 ,1107 ,2440 ,28229 ,27183 ,29807 ,9159 ,18085 ,15354 ,
      30684 ,5218 ,11609 ,954 ,24260 ,6069 ,23285 ,23363 ,1428 ,31086 ,28305 ,15273 ,23987 ,12370 ,6623 ,21065 ,29083 ,13194 ,6869 ,4009 ,27464 ,12014 ,31017 ,10792 ,32417 ,25762 ,17770 ,5534 ,29226 ,29964 ,27334 ,24569 ,7299 ,17125 ,18706 ,10385 ,9977 ,9663 ,6298 ,27740 ,32290 ,19558 ,17582 ,9714 ,27902 ,11964 ,1567 ,2996 ,32296 ,30279 ,13084 ,22124 ,25908 ,19917 ,8550 ,28787 ,15891 ,10309 ,23583 ,31587 ,16024 ,28256 ,18414 ,4086 ,18986 ,31954 ,28507 ,29490 ,22384 ,15967 ,14535 ,3159 ,7203 ,20684 ,854 ,12215 ,7977 ,11907 ,25870 ,21382 ,30215 ,14419 ,25471 ,13805 ,1721 ,27277 ,23514 ,17177 ,25622 ,12621 ,8735 ,8966 ,25358 ,21008 ,2793 ,13961 ,21445 ,27471 ,17490 ,15755 ,3681 ,12925 ,12409 ,28036 ,19899 ,11946 ,6051 ,29946 ,27259 ,11889 ,12907 ,12140 ,19564 ,7514 ,19346 ,13388 ,21259 ,8678 ,14500 ,19705 ,12982 ,22951 ,22318 ,9823 ,26633 ,12158 ,20090 ,28387 ,9021 ,22596 ,24874 ,18232 ,5972 ,22845 ,22693 ,30021 ,10092 ,23659 ,26815 ,11200 ,8152 ,12943 ,24787 ,20380 ,21720 ,9878 ,18524 ,23220 ,22019 ,3699 ,12071 ,5467 ,22760 ,16983 ,10772 ,19685 ,8414 ,32166 ,32203 ,1910 ,2516 ,23103 ,5589 ,28603 ,9343 ,12427 ,13939 ,21904 ,29541 ,18044 ,223 ,3823 ,16351 ,703 ,21564 ,10438 ,17588 ,2269 ,2975 ,31642 ,6126 ,26505 ,30913 ,17003 ,4303 ,26082 ,27925 ,2599 ,13546 ,28054 ,28656 ,16374 ,26823 ,7903 ,17952 ,28313 ,6587 ,17508 ,1183 ,25688 ,29927 ,8947 ,15254 ,31568 ,3804 ,19666 ,31549 ,14099 ,4388 ,6433 ,19974 ,16831 ,6921 ,14173 ,25289 ,22780 ,2911 ,25154 ,9252 ,6532 ,12643 ,15773 ,15455 ,27164 ,24166 ,12021 ,21284 ,18823 ,13657 ,14318 ,19740 ,1746 ,25933 ,6230 ,4756 ,14907 ,10918 ,27489 ,7382 ,31663 ,9720 ,30427 ,27002 ,6946 ,5869 ,21463 ,5894 ,2654 ,22233 ,22044 ,16073 ,14118 ,6151 ,1316 ,11088 ,7783 ,
      5599 ,31393 ,17682 ,24884 ,22490 ,17962 ,21294 ,26235 ,27632 ,28517 ,17500 ,4948 ,18716 ,8696 ,14230 ,11619 ,17918 ,18490 ,17456 ,13050 ,17483 ,21277 ,17439 ,17692 ,25228 ,5808 ,18463 ,17527 ,2732 ,26572 ,17709 ,15830 ,22301 ,14483 ,17473 ,12890 ,837 ,14518 ,25454 ,2776 ,17753 ,31000 ,11592 ,6606 ,17565 ,6281 ,13067 ,18397 ,27908 ,30896 ,5572 ,21547 ,26798 ,22676 ,18507 ,32186 ,9235 ,25272 ,17935 ,31532 ,4739 ,19723 ,26985 ,11071 ,32122 ,27676 ,18480 ,20210 ,18188 ,19364 ,8108 ,32070 ,23059 ,1844 ,21520 ,1202 ,16330 ,27238 ,17544 ,14688 ,14274 ,3211 ,4712 ,12756 ,14074 ,3455 ,5825 ,8434 ,25110 ,25132 ,25245 ,1373 ,25644 ,13406 ,29883 ,18760 ,11845 ,31024 ,17446 ,22534 ,13344 ,5746 ,26589 ,7105 ,14375 ,13320 ,2749 ,29160 ,21338 ,7532 ,18942 ,2290 ,11970 ,3578 ,17726 ,28915 ,15229 ,19582 ,24216 ,4162 ,19514 ,27546 ,6254 ,25707 ,28743 ,5643 ,15847 ,18068 ,11297 ,22854 ,17517 ,14026 ,15976 ,22336 ,3756 ,6078 ,19373 ,24375 ,1175 ,17971 ,29759 ,22345 ,4965 ,10699 ,27596 ,7167 ,18161 ,881 ,6408 ,30136 ,28534 ,32223 ,28824 ,8762 ,27649 ,12852 ,25498 ,9841 ,9410 ,23441 ,13111 ,16236 ,25218 ,8361 ,22902 ,23610 ,8713 ,13271 ,20594 ,29136 ,18733 ,30823 ,26482 ,22969 ,20431 ,17609 ,1573 ,17797 ,14247 ,12779 ,6896 ,13000 ,28134 ,20521 ,21773 ,13828 ,3428 ,28332 ,16854 ,10521 ,11636 ,9552 ,11208 ,29292 ,26562 ,15281 ,11503 ,4956 ,17979 ,370 ,6832 ,9279 ,22507 ,20792 ,20001 ,12176 ,9625 ,24469 ,15075 ,32502 ,21311 ,28111 ,6507 ,26651 ,21651 ,4783 ,27029 ,8853 ,13293 ,7922 ,11345 ,16100 ,26252 ,21926 ,12484 ,10799 ,17699 ,16633 ,18551 ,20108 ,31315 ,16905 ,3079 ,18918 ,4135 ,26842 ,14709 ,16752 ,24901 ,24066 ,3002 ,760 ,19487 ,13469 ,15430 ,27952 ,31410 ,1930 ,8040 ,19195 ,5616 ,20953 ,5062 ,28405 ,1063 ,250 ,
      29553 ,21133 ,18750 ,2528 ,29398 ,17600 ,4315 ,634 ,7012 ,21732 ,22772 ,4775 ,10104 ,7343 ,30840 ,9033 ,5693 ,4400 ,2923 ,10021 ,29939 ,14900 ,29153 ,26835 ,25945 ,20480 ,20611 ,24178 ,6342 ,9732 ,22245 ,18306 ,1611 ,30227 ,25634 ,15702 ,7215 ,32366 ,22986 ,18998 ,19911 ,8672 ,26499 ,21457 ,22670 ,19576 ,12994 ,27946 ,32302 ,32334 ,20448 ,7311 ,32392 ,32308 ,15903 ,3391 ,4602 ,29095 ,32429 ,14926 ,1440 ,576 ,17626 ,30696 ,30395 ,14286 ,25122 ,19634 ,23071 ,26473 ,23627 ,32134 ,14387 ,15935 ,22919 ,11857 ,5186 ,11982 ,19526 ,28224 ,17765 ,23578 ,8730 ,22313 ,10767 ,27920 ,9247 ,16068 ,18458 ,17930 ,25240 ,6249 ,27644 ,3423 ,13288 ,5611 ,20606 ,32424 ,25235 ,13123 ,8594 ,1585 ,21785 ,11687 ,31770 ,27608 ,28836 ,25952 ,19385 ,10618 ,8378 ,11309 ,30285 ,15087 ,27041 ,18635 ,6844 ,32340 ,16253 ,11220 ,3091 ,30095 ,13128 ,12496 ,23885 ,3014 ,8052 ,9127 ,16600 ,20759 ,12746 ,12819 ,20177 ,29127 ,13017 ,31499 ,28570 ,11167 ,6913 ,6499 ,921 ,9681 ,13772 ,9790 ,15176 ,4634 ,28151 ,17847 ,31061 ,9995 ,23812 ,2202 ,14821 ,24428 ,8599 ,27508 ,26308 ,13509 ,20538 ,4868 ,17311 ,28955 ,14264 ,19293 ,26731 ,6316 ,31932 ,29270 ,27378 ,26211 ,31139 ,10937 ,18209 ,14958 ,12796 ,24957 ,13090 ,11824 ,7278 ,24145 ,23962 ,20454 ,17814 ,23679 ,31868 ,32461 ,1590 ,23712 ,4458 ,27758 ,1119 ,21587 ,8160 ,1472 ,3445 ,23995 ,24533 ,18724 ,29767 ,22164 ,4049 ,5021 ,2015 ,7401 ,32736 ,7744 ,28349 ,15554 ,6667 ,14587 ,15519 ,11274 ,929 ,608 ,13845 ,10112 ,9466 ,13428 ,21790 ,24707 ,21030 ,10403 ,14653 ,24031 ,23733 ,25769 ,5815 ,24304 ,27080 ,6986 ,10538 ,12290 ,32036 ,17658 ,16871 ,20487 ,23329 ,17143 ,21870 ,2620 ,22130 ,2168 ,11653 ,3357 ,23260 ,7317 ,13707 ,2114 ,21191 ,16711 ,11692 ,31682 ,19092 ,30728 ,9569 ,488 ,
      6770 ,29697 ,32060 ,22428 ,2849 ,8352 ,30153 ,27402 ,31794 ,23018 ,6425 ,32494 ,14579 ,19935 ,17069 ,4216 ,32017 ,9447 ,28551 ,31849 ,19892 ,25926 ,14368 ,3072 ,31763 ,32029 ,31775 ,14337 ,31806 ,19030 ,32240 ,6782 ,31837 ,7247 ,18178 ,31901 ,15145 ,8568 ,20146 ,13741 ,32005 ,5784 ,19061 ,13676 ,8129 ,1984 ,898 ,14622 ,25914 ,2892 ,10073 ,4284 ,32271 ,32398 ,7184 ,12963 ,14356 ,25091 ,27613 ,9216 ,20575 ,28805 ,6813 ,8021 ,27390 ,17241 ,27666 ,17323 ,19272 ,13102 ,31880 ,25402 ,2837 ,15188 ,14833 ,19759 ,28582 ,15734 ,12869 ,16612 ,29685 ,6679 ,9478 ,10676 ,4061 ,9101 ,8779 ,8172 ,32048 ,25666 ,28841 ,23745 ,25380 ,22142 ,21203 ,26391 ,32482 ,17777 ,18470 ,3558 ,14399 ,30259 ,9858 ,30407 ,31782 ,2708 ,25515 ,20618 ,11438 ,30297 ,3103 ,26103 ,19923 ,1643 ,9427 ,1623 ,23558 ,32314 ,4614 ,2148 ,17057 ,5705 ,25957 ,1765 ,7024 ,31212 ,23458 ,29565 ,14610 ,22702 ,1192 ,4491 ,14544 ,23601 ,5151 ,23294 ,8117 ,27867 ,19966 ,21303 ,15511 ,3765 ,17988 ,6702 ,5772 ,12585 ,20829 ,3274 ,17100 ,19608 ,24392 ,24807 ,19049 ,11030 ,19390 ,7067 ,3314 ,31605 ,4247 ,3481 ,31889 ,29025 ,23049 ,30162 ,26168 ,5160 ,22362 ,11481 ,31825 ,13026 ,29776 ,27791 ,23636 ,10327 ,11144 ,4324 ,8556 ,1663 ,4982 ,3234 ,9952 ,15909 ,32525 ,26677 ,20134 ,14442 ,10623 ,18842 ,6456 ,27978 ,10716 ,7438 ,12951 ,19315 ,27228 ,12378 ,30184 ,8704 ,22353 ,25839 ,32259 ,18675 ,15993 ,8519 ,30653 ,28274 ,27433 ,27303 ,2880 ,19943 ,3773 ,1152 ,9689 ,16042 ,13626 ,7351 ,10061 ,24843 ,8383 ,12040 ,2485 ,192 ,6095 ,28625 ,9204 ,5541 ,17534 ,25423 ,17887 ,18432 ,22459 ,14199 ,14344 ,17415 ,28712 ,24185 ,32091 ,21489 ,14043 ,29852 ,28793 ,18130 ,29728 ,3725 ,1542 ,3397 ,22871 ,20400 ,6801 ,26531 ,11314 ,21620 ,12453 ,4104 ,15399 ,1032 ,
      7426 ,23114 ,2280 ,24636 ,9889 ,20512 ,26668 ,22607 ,6444 ,25581 ,6524 ,7914 ,24699 ,12032 ,30438 ,10962 ,14430 ,25977 ,21668 ,31965 ,11882 ,27482 ,7525 ,16745 ,10611 ,17136 ,30290 ,21482 ,13205 ,16448 ,4800 ,5229 ,3222 ,3957 ,21328 ,27687 ,32640 ,31035 ,3589 ,27816 ,8544 ,14494 ,30907 ,5888 ,18501 ,24210 ,28128 ,31404 ,15897 ,16247 ,17808 ,13701 ,7178 ,4608 ,32519 ,22865 ,32513 ,20643 ,15092 ,29303 ,19784 ,10810 ,771 ,10200 ,11469 ,6374 ,13310 ,26764 ,5938 ,6887 ,9943 ,21225 ,26156 ,3640 ,30328 ,5913 ,30505 ,16944 ,7939 ,13880 ,29013 ,12562 ,2363 ,7144 ,3134 ,9764 ,8870 ,5992 ,23037 ,29905 ,27046 ,23928 ,2815 ,4027 ,26134 ,1508 ,27779 ,29233 ,2739 ,15016 ,2397 ,16574 ,16117 ,19428 ,31813 ,22277 ,11362 ,6349 ,4526 ,13212 ,23184 ,28075 ,10315 ,1785 ,26269 ,25051 ,28482 ,29101 ,20649 ,6195 ,11132 ,8637 ,18640 ,2673 ,25546 ,18338 ,21943 ,26926 ,6690 ,11765 ,22524 ,17252 ,2343 ,17788 ,1654 ,12687 ,15499 ,7258 ,2903 ,27021 ,9458 ,10053 ,20809 ,29708 ,27855 ,29036 ,1674 ,19852 ,12596 ,24119 ,9296 ,22713 ,19954 ,2955 ,6849 ,19326 ,4692 ,5552 ,18141 ,19467 ,4479 ,28966 ,11835 ,8497 ,4645 ,4432 ,12193 ,20770 ,14598 ,18373 ,20018 ,1483 ,5444 ,25780 ,2179 ,13567 ,23589 ,5725 ,9642 ,14297 ,25333 ,32435 ,15098 ,31716 ,5139 ,30238 ,32345 ,6965 ,4411 ,16553 ,24486 ,21144 ,24795 ,28977 ,5736 ,6631 ,29047 ,14238 ,4973 ,11776 ,17088 ,29185 ,11520 ,28988 ,1227 ,29982 ,29452 ,5296 ,12573 ,17077 ,17996 ,6385 ,13780 ,29244 ,1796 ,30848 ,20817 ,3968 ,16258 ,30446 ,25988 ,26867 ,387 ,23125 ,7055 ,29971 ,26579 ,17344 ,12240 ,27352 ,5355 ,11726 ,19037 ,11568 ,31243 ,9739 ,20231 ,16455 ,15298 ,10147 ,31593 ,29441 ,12707 ,8312 ,23489 ,14932 ,29309 ,30041 ,4235 ,12329 ,11225 ,15653 ,8263 ,24587 ,29596 ,3848 ,
      28613 ,10136 ,4152 ,18242 ,2226 ,28323 ,18833 ,19126 ,2473 ,29500 ,15765 ,16092 ,10395 ,184 ,26859 ,964 ,24831 ,20220 ,22544 ,29645 ,12900 ,7375 ,18935 ,24894 ,8371 ,21863 ,3096 ,14036 ,23177 ,15291 ,16643 ,8196 ,1140 ,11557 ,15219 ,6016 ,8904 ,24507 ,16769 ,5405 ,2868 ,30872 ,14726 ,14991 ,22737 ,31104 ,14798 ,28677 ,16030 ,31232 ,24918 ,26351 ,21420 ,1446 ,19790 ,30786 ,13614 ,26041 ,30100 ,14137 ,14864 ,9065 ,24083 ,2052 ,25827 ,17333 ,3568 ,5334 ,31911 ,21764 ,20125 ,22438 ,30172 ,21978 ,18568 ,4501 ,13918 ,12388 ,25433 ,31294 ,19303 ,7044 ,31332 ,12829 ,12115 ,24005 ,24314 ,30762 ,27216 ,19644 ,13133 ,22063 ,15712 ,7722 ,16922 ,2538 ,8507 ,27341 ,17716 ,17262 ,10266 ,6641 ,17354 ,8458 ,32247 ,26774 ,15026 ,22252 ,27697 ,4807 ,16650 ,24646 ,28262 ,5344 ,17272 ,17201 ,6026 ,582 ,10816 ,18252 ,27421 ,22804 ,12501 ,24990 ,5491 ,21083 ,3907 ,15592 ,29840 ,30030 ,25697 ,24980 ,3168 ,10512 ,27969 ,23372 ,32079 ,4347 ,15447 ,26244 ,14645 ,6087 ,379 ,30585 ,17403 ,23478 ,31427 ,11398 ,7489 ,24278 ,23776 ,13590 ,28700 ,27123 ,23890 ,1335 ,28872 ,666 ,1947 ,20283 ,25411 ,29430 ,19504 ,27411 ,30957 ,23303 ,25848 ,9603 ,9192 ,31508 ,22173 ,6170 ,32143 ,20320 ,13486 ,643 ,18420 ,12696 ,11785 ,3518 ,21234 ,17632 ,777 ,22616 ,22447 ,7862 ,3019 ,19135 ,4905 ,23381 ,26422 ,10461 ,20388 ,15642 ,5633 ,21073 ,16193 ,11627 ,10707 ,26413 ,1530 ,10877 ,14761 ,11107 ,9509 ,2560 ,20970 ,7684 ,18118 ,4224 ,6710 ,9387 ,9798 ,2088 ,19212 ,9041 ,29716 ,18782 ,8057 ,10970 ,13983 ,972 ,30593 ,132 ,21608 ,24576 ,15837 ,3897 ,8810 ,21165 ,28422 ,16514 ,6789 ,26961 ,5079 ,18313 ,327 ,5236 ,8203 ,16395 ,4092 ,29585 ,1080 ,31172 ,20065 ,30702 ,10206 ,522 ,15387 ,1275 ,9132 ,7802 ,20910 ,72 ,267 ,12 ,
      15342 ,477 ,28377 ,26916 ,16148 ,11062 ,8012 ,2043 ,29795 ,30540 ,1902 ,23433 ,4860 ,3473 ,19459 ,20275 ,2428 ,19081 ,18890 ,21818 ,21375 ,14092 ,14681 ,24462 ,28217 ,15547 ,16605 ,27296 ,13873 ,5289 ,31287 ,7677 ,10566 ,16700 ,26623 ,25536 ,32595 ,5843 ,15047 ,4563 ,27734 ,28030 ,21898 ,1740 ,2770 ,7099 ,13265 ,16899 ,18992 ,11681 ,29264 ,12284 ,13735 ,30401 ,11475 ,14193 ,27810 ,19422 ,20764 ,11720 ,5399 ,8452 ,9597 ,16508 ,4557 ,3346 ,22941 ,8627 ,29353 ,4730 ,20566 ,14855 ,30350 ,28179 ,13243 ,23533 ,23840 ,18590 ,25190 ,10573 ,4004 ,22119 ,13800 ,13383 ,23215 ,31637 ,16826 ,6941 ,13045 ,21542 ,12751 ,28910 ,876 ,12774 ,28106 ,13464 ,10016 ,7306 ,22308 ,18630 ,17842 ,24140 ,11269 ,3352 ,31844 ,4279 ,10671 ,1618 ,3269 ,3229 ,1147 ,3720 ,31960 ,13696 ,7139 ,25046 ,19847 ,14292 ,6380 ,8307 ,29640 ,26346 ,12824 ,17196 ,11393 ,3513 ,9382 ,31167 ,21813 ,12279 ,13378 ,25041 ,7585 ,25263 ,25082 ,26032 ,431 ,7631 ,8406 ,25490 ,26300 ,3306 ,4684 ,28864 ,32679 ,27069 ,1816 ,7590 ,16281 ,16805 ,16302 ,25309 ,10346 ,20861 ,20182 ,13156 ,32687 ,1391 ,8080 ,2436 ,31082 ,25758 ,19554 ,10305 ,20680 ,12617 ,11942 ,22947 ,23655 ,16979 ,18040 ,26078 ,8943 ,25150 ,6226 ,22040 ,28513 ,5804 ,30996 ,25268 ,1840 ,25128 ,13316 ,27542 ,24371 ,8758 ,29132 ,13824 ,9275 ,8849 ,18914 ,19191 ,21728 ,20476 ,8668 ,29091 ,15931 ,17926 ,27604 ,30091 ,11163 ,24424 ,26207 ,32457 ,5017 ,13424 ,17654 ,16707 ,23014 ,32025 ,5780 ,25087 ,15184 ,25662 ,2704 ,5701 ,27863 ,11026 ,13022 ,14438 ,18671 ,24839 ,17411 ,26527 ,25577 ,17132 ,14490 ,20639 ,3636 ,29901 ,22273 ,8633 ,7254 ,2951 ,18369 ,30234 ,29181 ,3964 ,11564 ,12325 ,29496 ,21859 ,30868 ,26037 ,21974 ,19640 ,26770 ,22800 ,4343 ,27119 ,31504 ,7858 ,10873 ,18778 ,26957 ,1271 ,
      30536 ,15543 ,28026 ,19418 ,28175 ,21538 ,4275 ,26342 ,7627 ,20857 ,16975 ,8754 ,24420 ,11022 ,2947 ,27115 ,20853 ,32725 ,18016 ,436 ,7970 ,3797 ,16323 ,19994 ,5179 ,32729 ,28575 ,30646 ,30498 ,1220 ,13911 ,9502 ,23833 ,5010 ,3671 ,2387 ,32553 ,9317 ,21692 ,29359 ,26187 ,18020 ,1882 ,10651 ,1698 ,1862 ,10744 ,12092 ,22390 ,2004 ,22568 ,7636 ,20722 ,23077 ,5944 ,31356 ,31451 ,440 ,11172 ,8985 ,30359 ,6734 ,24759 ,29804 ,24257 ,23984 ,27461 ,29223 ,9974 ,27899 ,25905 ,16021 ,22381 ,7974 ,1718 ,25355 ,3678 ,27256 ,21256 ,26630 ,5969 ,8149 ,22016 ,8411 ,9340 ,16348 ,6123 ,13543 ,6584 ,3801 ,6918 ,12640 ,13654 ,10915 ,5866 ,6148 ,22487 ,18713 ,17480 ,2729 ,834 ,17562 ,26795 ,4736 ,18185 ,16327 ,14071 ,25641 ,13341 ,21335 ,15226 ,28740 ,15973 ,29756 ,6405 ,25495 ,22899 ,26479 ,6893 ,16851 ,11500 ,19998 ,6504 ,11342 ,18548 ,14706 ,15427 ,5059 ,29395 ,10101 ,29936 ,6339 ,7212 ,22667 ,32389 ,1437 ,23068 ,5183 ,10764 ,27641 ,8591 ,19382 ,6841 ,23882 ,20174 ,918 ,31058 ,26305 ,26728 ,18206 ,23959 ,4455 ,24530 ,32733 ,926 ,21027 ,27077 ,23326 ,23257 ,19089 ,2846 ,14576 ,19889 ,31803 ,15142 ,8126 ,32268 ,20572 ,19269 ,28579 ,4058 ,25377 ,14396 ,11435 ,23555 ,7021 ,14541 ,15508 ,17097 ,3311 ,26165 ,23633 ,9949 ,6453 ,30181 ,30650 ,9686 ,2482 ,17884 ,32088 ,1539 ,12450 ,9886 ,24696 ,11879 ,13202 ,32637 ,18498 ,7175 ,19781 ,5935 ,30502 ,3131 ,2812 ,2394 ,4523 ,28479 ,25543 ,2340 ,9455 ,12593 ,4689 ,4642 ,5441 ,25330 ,4408 ,29044 ,1224 ,13777 ,25985 ,12237 ,20228 ,23486 ,8260 ,2223 ,10392 ,12897 ,23174 ,8901 ,22734 ,21417 ,14861 ,31908 ,13915 ,12112 ,15709 ,10263 ,27694 ,6023 ,5488 ,3165 ,14642 ,7486 ,28869 ,30954 ,32140 ,21231 ,4902 ,16190 ,9506 ,9795 ,13980 ,8807 ,324 ,20062 ,20907 ,
      16145 ,4857 ,21372 ,13870 ,32592 ,2767 ,13732 ,5396 ,29350 ,23837 ,23212 ,873 ,17839 ,3266 ,19844 ,11390 ,7582 ,26297 ,16278 ,32684 ,20677 ,8940 ,1837 ,9272 ,15928 ,5014 ,15181 ,18668 ,3633 ,29178 ,21971 ,10870 ,28172 ,24417 ,7967 ,30495 ,32550 ,1695 ,20719 ,30356 ,9971 ,3675 ,9337 ,13651 ,831 ,13338 ,22896 ,18545 ,7209 ,8588 ,26725 ,27074 ,15139 ,14393 ,26162 ,17881 ,32634 ,2391 ,4639 ,12234 ,8898 ,10260 ,30951 ,8804 ,32589 ,17836 ,20674 ,3630 ,32547 ,828 ,15136 ,8895 ,32544 ,32557 ,32573 ,15120 ,32560 ,7550 ,799 ,32602 ,3617 ,15165 ,7566 ,1821 ,32576 ,21356 ,29334 ,19828 ,815 ,9321 ,28156 ,20703 ,15123 ,26709 ,32618 ,30935 ,19815 ,9984 ,844 ,30318 ,32563 ,18960 ,4828 ,28185 ,15152 ,21696 ,10841 ,7222 ,7553 ,32647 ,8911 ,24339 ,20690 ,23801 ,30466 ,7595 ,802 ,15941 ,3646 ,6552 ,26696 ,29363 ,17852 ,19237 ,32605 ,2308 ,10231 ,16158 ,10857 ,31488 ,29480 ,26754 ,3620 ,14474 ,7238 ,11548 ,5001 ,26191 ,21712 ,27588 ,15168 ,5764 ,27847 ,17395 ,32671 ,20166 ,32663 ,16286 ,7569 ,13362 ,415 ,4668 ,8927 ,18024 ,31066 ,11926 ,1824 ,30980 ,24355 ,18898 ,5383 ,20748 ,18976 ,11459 ,32579 ,26607 ,27718 ,13249 ,4844 ,1886 ,15326 ,7996 ,21359 ,18874 ,28201 ,31271 ,860 ,12735 ,3988 ,16810 ,29337 ,22925 ,30334 ,25174 ,3253 ,10655 ,10000 ,11253 ,19831 ,7123 ,29624 ,9366 ,18532 ,6488 ,15957 ,6877 ,818 ,17464 ,18169 ,15210 ,3662 ,1702 ,24241 ,25889 ,9324 ,22000 ,6568 ,5850 ,30482 ,28559 ,20837 ,16307 ,28159 ,28010 ,7611 ,2931 ,1682 ,1866 ,23817 ,21676 ,20706 ,22552 ,31435 ,24743 ,17868 ,9670 ,14525 ,9933 ,15126 ,19873 ,19253 ,23539 ,8575 ,10748 ,29379 ,32373 ,26712 ,31042 ,24514 ,23241 ,12221 ,13761 ,2324 ,25314 ,32621 ,11863 ,5919 ,28463 ,10247 ,12096 ,2207 ,21401 ,30938 ,7470 ,16174 ,20046 ,
      9353 ,24946 ,17167 ,5982 ,19818 ,6597 ,13667 ,14982 ,10642 ,22394 ,3691 ,30128 ,9987 ,19600 ,24111 ,24270 ,16797 ,18198 ,13354 ,10351 ,847 ,15247 ,21513 ,22500 ,22912 ,2008 ,14826 ,15986 ,30321 ,11513 ,18561 ,14754 ,13236 ,26200 ,1711 ,3124 ,32566 ,24234 ,16671 ,23846 ,20735 ,22572 ,16479 ,22403 ,18963 ,31464 ,30372 ,25804 ,7983 ,31128 ,26887 ,20866 ,4831 ,5192 ,30511 ,15793 ,18861 ,7640 ,24433 ,20344 ,28188 ,4180 ,5260 ,30549 ,17382 ,19282 ,14409 ,12552 ,15155 ,17744 ,31996 ,2859 ,26178 ,20726 ,16678 ,14554 ,21699 ,30194 ,17897 ,15054 ,26741 ,17300 ,26008 ,20187 ,10844 ,24543 ,27090 ,12663 ,14461 ,23081 ,8604 ,12529 ,7225 ,28933 ,3935 ,29408 ,4655 ,6305 ,25461 ,2353 ,7556 ,29057 ,12250 ,18596 ,20153 ,5948 ,2407 ,22993 ,32650 ,3596 ,16776 ,9899 ,11913 ,31921 ,10276 ,13161 ,8914 ,11988 ,16950 ,2236 ,30967 ,31360 ,27513 ,3178 ,24342 ,16203 ,8820 ,727 ,24730 ,23668 ,8956 ,23918 ,20693 ,6272 ,1975 ,31095 ,1853 ,31455 ,12063 ,28526 ,23804 ,24384 ,9288 ,23768 ,16294 ,23951 ,407 ,32692 ,30469 ,10359 ,32700 ,15475 ,27997 ,444 ,26313 ,22086 ,7598 ,25725 ,10993 ,21826 ,15197 ,11813 ,25612 ,23027 ,805 ,27876 ,18684 ,25196 ,6475 ,11176 ,5030 ,3047 ,15944 ,27564 ,26450 ,21741 ,25876 ,7267 ,29194 ,1396 ,3649 ,19532 ,7945 ,25590 ,21987 ,8989 ,13514 ,29509 ,6555 ,4356 ,10886 ,22201 ,23228 ,23701 ,20998 ,4017 ,26699 ,13058 ,889 ,14789 ,10735 ,30363 ,23853 ,31738 ,29366 ,5661 ,22638 ,4570 ,9920 ,31857 ,3282 ,8085 ,17855 ,28761 ,30621 ,10029 ,19860 ,6738 ,20543 ,31973 ,19240 ,29653 ,11406 ,17025 ,28450 ,27747 ,2783 ,26124 ,32608 ,15865 ,24667 ,10579 ,13748 ,24763 ,8231 ,19005 ,2311 ,27823 ,5412 ,5107 ,21388 ,1108 ,23145 ,2441 ,10234 ,28230 ,13886 ,27184 ,7457 ,29808 ,4873 ,9160 ,16161 ,18086 ,295 ,15355 ,
      1258 ,30685 ,24559 ,5219 ,10860 ,11610 ,4207 ,955 ,27106 ,24261 ,30013 ,6070 ,31491 ,23286 ,12679 ,23364 ,26024 ,1429 ,11540 ,31087 ,29483 ,28306 ,20203 ,15274 ,19627 ,23988 ,17316 ,12371 ,26757 ,6624 ,5327 ,21066 ,8620 ,29084 ,29216 ,13195 ,3623 ,6870 ,12545 ,4010 ,17119 ,27465 ,23097 ,12015 ,14477 ,31018 ,16230 ,10793 ,30221 ,32418 ,28949 ,25763 ,7241 ,17771 ,29019 ,5535 ,3951 ,29227 ,28960 ,29965 ,11551 ,27335 ,29424 ,24570 ,16694 ,7300 ,25752 ,17126 ,5004 ,18707 ,14570 ,10386 ,24411 ,9978 ,20742 ,9664 ,26194 ,6299 ,11807 ,27741 ,29078 ,32291 ,30210 ,19559 ,21715 ,17583 ,4383 ,9715 ,17913 ,27903 ,14269 ,11965 ,27591 ,1568 ,15070 ,2997 ,5688 ,32297 ,17760 ,30280 ,15171 ,13085 ,6662 ,22125 ,32012 ,25909 ,29680 ,19918 ,5767 ,8551 ,2875 ,28788 ,14425 ,15892 ,29008 ,10310 ,27850 ,23584 ,12568 ,31588 ,24826 ,16025 ,19298 ,28257 ,17398 ,18415 ,18113 ,4087 ,2423 ,18987 ,3999 ,31955 ,32674 ,28508 ,23009 ,29491 ,20848 ,22385 ,5964 ,15968 ,20169 ,14536 ,2335 ,3160 ,7577 ,7204 ,3612 ,20685 ,32666 ,855 ,30477 ,12216 ,16792 ,7978 ,26736 ,11908 ,16289 ,25871 ,9915 ,21383 ,26019 ,30216 ,29073 ,14420 ,7572 ,25472 ,10287 ,13806 ,12266 ,1722 ,26898 ,27278 ,13365 ,23515 ,18612 ,17178 ,25477 ,25623 ,29205 ,12622 ,418 ,8736 ,2369 ,8967 ,3293 ,25359 ,6321 ,21009 ,4671 ,2794 ,23156 ,13962 ,22027 ,21446 ,12004 ,27472 ,8930 ,17491 ,6416 ,15756 ,16966 ,3682 ,22579 ,12926 ,18027 ,12410 ,2252 ,28037 ,10292 ,19900 ,17108 ,11947 ,31069 ,6052 ,13177 ,29947 ,12604 ,27260 ,31937 ,11890 ,11929 ,12908 ,7497 ,12141 ,27529 ,19565 ,31007 ,7515 ,1827 ,19347 ,3194 ,13389 ,5791 ,21260 ,31376 ,8679 ,30983 ,14501 ,30879 ,19706 ,13811 ,12983 ,16219 ,22952 ,24358 ,22319 ,7150 ,9824 ,8836 ,26634 ,29275 ,12159 ,18901 ,20091 ,743 ,28388 ,
      16495 ,9022 ,23353 ,22597 ,5386 ,24875 ,22419 ,18233 ,19409 ,5973 ,22588 ,22846 ,20751 ,22694 ,11757 ,30022 ,12271 ,10093 ,31480 ,23660 ,18979 ,26816 ,32115 ,11201 ,30388 ,8153 ,27383 ,12944 ,11462 ,24788 ,25820 ,20381 ,4550 ,21721 ,24250 ,9879 ,32582 ,18525 ,17375 ,23221 ,16687 ,22020 ,20255 ,3700 ,26610 ,12072 ,23862 ,5468 ,1727 ,22761 ,30002 ,16984 ,27721 ,10773 ,3140 ,19686 ,7086 ,8415 ,26216 ,32167 ,13252 ,32204 ,351 ,1911 ,20262 ,2517 ,5208 ,23104 ,4847 ,5590 ,6761 ,28604 ,30527 ,9344 ,16486 ,12428 ,1889 ,13940 ,15809 ,21905 ,26903 ,29542 ,1247 ,18045 ,15329 ,224 ,20882 ,3824 ,11049 ,16352 ,31144 ,704 ,7999 ,21565 ,10178 ,10439 ,24449 ,17589 ,11599 ,2270 ,21362 ,2976 ,20360 ,31643 ,19068 ,6127 ,7656 ,26506 ,18877 ,30914 ,14733 ,17004 ,27283 ,4304 ,4196 ,26083 ,28204 ,27926 ,9770 ,2600 ,5276 ,13547 ,10942 ,28055 ,31274 ,28657 ,30565 ,16375 ,13451 ,26824 ,15263 ,7904 ,863 ,17953 ,8343 ,28314 ,21529 ,6588 ,24866 ,17509 ,12738 ,1184 ,22516 ,25689 ,13370 ,29928 ,29472 ,8948 ,3991 ,15255 ,10367 ,31569 ,31624 ,3805 ,18214 ,19667 ,16813 ,31550 ,18805 ,14100 ,14842 ,4389 ,1418 ,6434 ,29340 ,19975 ,16002 ,16832 ,3333 ,6922 ,2024 ,14174 ,22928 ,25290 ,30072 ,22781 ,23520 ,2912 ,11529 ,25155 ,30337 ,9253 ,8876 ,6533 ,18577 ,12644 ,14963 ,15774 ,25177 ,15456 ,14770 ,27165 ,3707 ,24167 ,12360 ,12022 ,3256 ,21285 ,30144 ,18824 ,4266 ,13658 ,22410 ,14319 ,10658 ,19741 ,3540 ,1747 ,18617 ,25934 ,19616 ,6231 ,10003 ,4757 ,15684 ,14908 ,24127 ,10919 ,12801 ,27490 ,11256 ,7383 ,24286 ,31664 ,8294 ,9721 ,6613 ,30428 ,19834 ,27003 ,8479 ,6947 ,13683 ,5870 ,24618 ,21464 ,7126 ,5895 ,14998 ,2655 ,17183 ,22234 ,5316 ,22045 ,29627 ,16074 ,5998 ,14119 ,3500 ,6152 ,24962 ,1317 ,9369 ,11089 ,3879 ,7784 ,
      5046 ,5600 ,2986 ,31394 ,18535 ,17683 ,3063 ,24885 ,19985 ,22491 ,11192 ,17963 ,6491 ,21295 ,27013 ,26236 ,25482 ,27633 ,27580 ,28518 ,15960 ,17501 ,19357 ,4949 ,26466 ,18717 ,13095 ,8697 ,6880 ,14231 ,21757 ,11620 ,4723 ,17919 ,27892 ,18491 ,821 ,17457 ,17737 ,13051 ,18700 ,17484 ,5583 ,21278 ,17467 ,17440 ,25212 ,17693 ,25628 ,25229 ,14258 ,5809 ,18172 ,18464 ,23043 ,17528 ,21322 ,2733 ,11829 ,26573 ,15213 ,17710 ,19498 ,15831 ,26617 ,22302 ,19548 ,14484 ,3665 ,17474 ,19883 ,12891 ,7961 ,838 ,18970 ,14519 ,1705 ,25455 ,25606 ,2777 ,29210 ,17754 ,29067 ,31001 ,24244 ,11593 ,1412 ,6607 ,27886 ,17566 ,7283 ,6282 ,25892 ,13068 ,15875 ,18398 ,13530 ,27909 ,17572 ,30897 ,9327 ,5573 ,29525 ,21548 ,8136 ,26799 ,9005 ,22677 ,22003 ,18508 ,22744 ,32187 ,12627 ,9236 ,4372 ,25273 ,6571 ,17936 ,29911 ,31533 ,10902 ,4740 ,24150 ,19724 ,5853 ,26986 ,22217 ,11072 ,9489 ,32123 ,10375 ,27677 ,30485 ,18481 ,9438 ,20211 ,32716 ,18189 ,10084 ,19365 ,28562 ,8109 ,15491 ,32071 ,423 ,23060 ,4993 ,1845 ,20840 ,21521 ,32708 ,1203 ,3784 ,16331 ,23967 ,27239 ,16310 ,17545 ,29739 ,14689 ,26329 ,14275 ,7289 ,3212 ,28162 ,4713 ,22102 ,12757 ,15530 ,14075 ,460 ,3456 ,28013 ,5826 ,11664 ,8435 ,8741 ,25111 ,25741 ,25133 ,7614 ,25246 ,27052 ,1374 ,11009 ,25645 ,20459 ,13407 ,2934 ,29884 ,21842 ,18761 ,12079 ,11846 ,9653 ,31025 ,1685 ,17447 ,28542 ,22535 ,18007 ,13345 ,31471 ,5747 ,1869 ,26590 ,12718 ,7106 ,2374 ,14376 ,24400 ,13321 ,23820 ,2750 ,26280 ,29161 ,9304 ,21339 ,17819 ,7533 ,21679 ,18943 ,23784 ,2291 ,31343 ,11971 ,6288 ,3579 ,20709 ,17727 ,17283 ,28916 ,1991 ,15230 ,24929 ,19583 ,22555 ,24217 ,31111 ,4163 ,8972 ,19515 ,11796 ,27547 ,31438 ,6255 ,23934 ,25708 ,6721 ,28744 ,23684 ,5644 ,24746 ,15848 ,1091 ,18069 ,
      12437 ,11298 ,28777 ,22855 ,17871 ,17518 ,14328 ,14027 ,30637 ,15977 ,12935 ,22337 ,9673 ,3757 ,10045 ,6079 ,3298 ,19374 ,5756 ,24376 ,14528 ,1176 ,8101 ,17972 ,23620 ,29760 ,31873 ,22346 ,9936 ,4966 ,20118 ,10700 ,20559 ,27597 ,25898 ,7168 ,15129 ,18162 ,31989 ,882 ,14563 ,6409 ,6754 ,30137 ,19876 ,28535 ,31747 ,32224 ,25364 ,28825 ,29669 ,8763 ,19256 ,27650 ,2821 ,12853 ,11422 ,25499 ,32466 ,9842 ,23542 ,9411 ,17041 ,23442 ,23869 ,13112 ,30269 ,16237 ,8578 ,25219 ,31754 ,8362 ,5170 ,22903 ,30379 ,23611 ,10751 ,8714 ,18442 ,13272 ,6326 ,20595 ,5677 ,29137 ,29382 ,18734 ,6996 ,30824 ,22654 ,26483 ,1595 ,22970 ,32376 ,20432 ,4586 ,17610 ,4442 ,1574 ,13074 ,17798 ,26715 ,14248 ,27362 ,12780 ,905 ,6897 ,16584 ,13001 ,31045 ,28135 ,14805 ,20522 ,21014 ,21774 ,6651 ,13829 ,24517 ,3429 ,4033 ,28333 ,23313 ,16855 ,23717 ,10522 ,23244 ,11637 ,21175 ,9553 ,8247 ,11209 ,31577 ,29293 ,12224 ,26563 ,19021 ,15282 ,1211 ,11504 ,24779 ,4957 ,13764 ,17980 ,20801 ,371 ,4676 ,6833 ,27839 ,9280 ,2327 ,22508 ,15483 ,20793 ,5428 ,20002 ,4463 ,12177 ,25317 ,9626 ,5123 ,24470 ,19768 ,15076 ,15881 ,32503 ,32624 ,21312 ,8528 ,28112 ,24683 ,6508 ,7410 ,26652 ,11866 ,21652 ,10595 ,4784 ,2799 ,27030 ,28997 ,8854 ,5922 ,13294 ,26140 ,7923 ,4510 ,11346 ,27763 ,16101 ,28466 ,26253 ,11116 ,21927 ,5475 ,12485 ,28246 ,10800 ,10250 ,17700 ,32231 ,16634 ,13902 ,18552 ,25811 ,20109 ,12099 ,31316 ,27200 ,16906 ,23161 ,3080 ,24815 ,18919 ,2210 ,4136 ,2457 ,26843 ,22721 ,14710 ,1124 ,16753 ,21404 ,24902 ,13598 ,24067 ,4889 ,3003 ,18404 ,761 ,30941 ,19488 ,9176 ,13470 ,14629 ,15431 ,29824 ,27953 ,7473 ,31411 ,28684 ,1931 ,13967 ,8041 ,18102 ,19196 ,16177 ,5617 ,1514 ,20954 ,311 ,5063 ,21592 ,28406 ,20049 ,1064 ,15371 ,251 ,
      7771 ,29554 ,16364 ,21134 ,9356 ,18751 ,26382 ,2529 ,6139 ,29399 ,10430 ,17601 ,24949 ,4316 ,13559 ,635 ,22032 ,7013 ,31263 ,21733 ,17170 ,22773 ,8427 ,4776 ,16061 ,10105 ,8165 ,7344 ,5985 ,30841 ,30755 ,9034 ,6934 ,5694 ,13536 ,4401 ,19821 ,2924 ,12656 ,10022 ,9708 ,29940 ,3817 ,14901 ,6600 ,29154 ,30817 ,26836 ,21451 ,25946 ,10931 ,20481 ,13670 ,20612 ,27785 ,24179 ,5882 ,6343 ,1477 ,9733 ,14985 ,22246 ,6164 ,18307 ,1734 ,1612 ,26072 ,30228 ,10645 ,25635 ,25371 ,15703 ,13645 ,7216 ,7990 ,32367 ,22397 ,22987 ,3041 ,18999 ,12009 ,19912 ,27272 ,8673 ,3694 ,26500 ,14168 ,21458 ,21272 ,22671 ,3450 ,19577 ,30131 ,12995 ,26646 ,27947 ,14895 ,32303 ,27915 ,32335 ,9990 ,20449 ,603 ,7312 ,25921 ,32393 ,9096 ,32309 ,19603 ,15904 ,16037 ,3392 ,27477 ,4603 ,9759 ,29096 ,24114 ,32430 ,29239 ,14927 ,7370 ,1441 ,24000 ,577 ,24273 ,17627 ,2083 ,30697 ,14087 ,30396 ,31632 ,14287 ,16800 ,25123 ,25657 ,19635 ,3792 ,23072 ,16343 ,26474 ,18201 ,23628 ,5436 ,32135 ,8935 ,14388 ,21351 ,15936 ,13357 ,22920 ,28005 ,11858 ,15242 ,5187 ,24538 ,11983 ,10354 ,19527 ,28756 ,28225 ,28301 ,17766 ,17578 ,23579 ,850 ,8731 ,6047 ,22314 ,26811 ,10768 ,219 ,27921 ,15250 ,9248 ,4752 ,16069 ,17496 ,18459 ,11588 ,17931 ,21516 ,25241 ,2745 ,6250 ,1171 ,27645 ,18729 ,3424 ,22503 ,13289 ,4131 ,5612 ,22768 ,20607 ,26495 ,32425 ,22915 ,25236 ,28832 ,13124 ,6909 ,8595 ,31135 ,1586 ,2011 ,21786 ,16867 ,11688 ,6421 ,31771 ,19057 ,27609 ,14829 ,28837 ,25511 ,25953 ,19962 ,19386 ,29772 ,10619 ,15989 ,8379 ,28708 ,11310 ,6520 ,30286 ,30903 ,15088 ,30324 ,27042 ,11358 ,18636 ,2899 ,6845 ,20014 ,32341 ,11516 ,16254 ,31239 ,11221 ,15761 ,3092 ,14722 ,30096 ,18564 ,13129 ,15022 ,12497 ,15443 ,23886 ,22169 ,3015 ,14757 ,8053 ,5075 ,9128 ,
      1898 ,16601 ,21894 ,20760 ,13239 ,12747 ,10667 ,12820 ,8402 ,20178 ,18036 ,29128 ,26203 ,13018 ,18365 ,31500 ,16971 ,28571 ,1878 ,11168 ,1714 ,6914 ,14067 ,6500 ,10760 ,922 ,4054 ,9682 ,3127 ,13773 ,12108 ,9791 ,23208 ,15177 ,9333 ,4635 ,32569 ,28152 ,10837 ,17848 ,21708 ,31062 ,15322 ,9996 ,24237 ,23813 ,29375 ,2203 ,3687 ,14822 ,16475 ,24429 ,16674 ,8600 ,2403 ,27509 ,12059 ,26309 ,5026 ,13510 ,23849 ,20539 ,8227 ,4869 ,30009 ,17312 ,23093 ,28956 ,20738 ,14265 ,29676 ,19294 ,5960 ,26732 ,26894 ,6317 ,22575 ,31933 ,31372 ,29271 ,22584 ,27379 ,20251 ,26212 ,16482 ,31140 ,7652 ,10938 ,24862 ,18210 ,2020 ,14959 ,22406 ,12797 ,24614 ,24958 ,11188 ,13091 ,5579 ,11825 ,18966 ,7279 ,9001 ,24146 ,10080 ,23963 ,456 ,20455 ,31467 ,17815 ,24925 ,23680 ,12931 ,31869 ,6750 ,32462 ,30375 ,1591 ,16580 ,23713 ,24775 ,4459 ,7406 ,27759 ,25807 ,1120 ,29820 ,21588 ,10426 ,8161 ,3813 ,1473 ,7986 ,3446 ,9092 ,23996 ,16339 ,24534 ,215 ,18725 ,31131 ,29768 ,20010 ,22165 ,18032 ,4050 ,15318 ,5022 ,26890 ,2016 ,452 ,7402 ,211 ,32737 ,32741 ,7745 ,20869 ,28350 ,995 ,15555 ,28591 ,6668 ,29531 ,14588 ,4834 ,15520 ,30662 ,11275 ,2504 ,930 ,32745 ,609 ,5195 ,13846 ,21110 ,10113 ,12415 ,9467 ,1236 ,13429 ,30514 ,21791 ,16123 ,24708 ,13927 ,21031 ,7749 ,10404 ,15796 ,14654 ,9518 ,24032 ,16991 ,23734 ,693 ,25770 ,18864 ,5816 ,8770 ,24305 ,6114 ,27081 ,20873 ,6987 ,7643 ,10539 ,19157 ,12291 ,2257 ,32037 ,11038 ,17659 ,24436 ,16872 ,23408 ,20488 ,2963 ,23330 ,28354 ,17144 ,20347 ,21871 ,27131 ,2621 ,2587 ,22131 ,21554 ,2169 ,28191 ,11654 ,18273 ,3358 ,4291 ,23261 ,999 ,7318 ,4183 ,13708 ,26358 ,2115 ,28042 ,21192 ,10167 ,16712 ,5263 ,11693 ,19434 ,31683 ,28644 ,19093 ,15559 ,30729 ,30552 ,9570 ,99 ,489 ,
      4074 ,6771 ,20370 ,29698 ,17385 ,32061 ,25393 ,22429 ,16012 ,2850 ,28595 ,8353 ,19285 ,30154 ,8489 ,27403 ,10297 ,31795 ,11451 ,23019 ,14412 ,6426 ,3204 ,32495 ,23571 ,14580 ,6672 ,19936 ,12555 ,17070 ,7037 ,4217 ,22112 ,32018 ,8142 ,9448 ,15158 ,28552 ,17293 ,31850 ,32284 ,19893 ,29535 ,25927 ,17747 ,14369 ,20588 ,3073 ,19905 ,31764 ,27372 ,32030 ,31999 ,31776 ,31819 ,14338 ,8538 ,31807 ,14592 ,19031 ,2862 ,32241 ,9186 ,6783 ,27728 ,31838 ,23649 ,7248 ,26181 ,18179 ,19263 ,31902 ,9965 ,15146 ,4838 ,8569 ,20729 ,20147 ,6469 ,13742 ,17113 ,32006 ,12260 ,5785 ,16681 ,19062 ,3327 ,13677 ,18694 ,8130 ,15524 ,1985 ,14557 ,899 ,24677 ,14623 ,9702 ,25915 ,26805 ,2893 ,21702 ,10074 ,2498 ,4285 ,32278 ,32272 ,30666 ,32399 ,30197 ,7185 ,21427 ,12964 ,11952 ,14357 ,32104 ,25092 ,17900 ,27614 ,22283 ,9217 ,1555 ,20576 ,11279 ,28806 ,15057 ,6814 ,12466 ,8022 ,21053 ,27391 ,18222 ,17242 ,26744 ,27667 ,17232 ,17324 ,23975 ,19273 ,2508 ,13103 ,17303 ,31881 ,4471 ,25403 ,31074 ,2838 ,5375 ,15189 ,26011 ,14834 ,26321 ,19760 ,28293 ,28583 ,934 ,15735 ,20190 ,12870 ,14006 ,16613 ,942 ,29686 ,9011 ,6680 ,10847 ,9479 ,21043 ,10677 ,30672 ,4062 ,32749 ,9102 ,24546 ,8780 ,18283 ,8173 ,6057 ,32049 ,23342 ,25667 ,27093 ,28842 ,11368 ,23746 ,23273 ,25381 ,613 ,22143 ,12666 ,21204 ,19105 ,26392 ,10780 ,32483 ,22835 ,17778 ,14464 ,18471 ,27657 ,3559 ,27452 ,14400 ,5199 ,30260 ,23084 ,9859 ,7884 ,30408 ,13182 ,31783 ,19398 ,2709 ,8607 ,25516 ,25021 ,20619 ,6857 ,11439 ,13850 ,30298 ,12532 ,3104 ,23898 ,26104 ,5522 ,19924 ,22683 ,1644 ,7228 ,9428 ,17222 ,1624 ,32405 ,23559 ,21114 ,32315 ,28936 ,4615 ,1453 ,2149 ,29952 ,17058 ,11746 ,5706 ,3938 ,25958 ,6355 ,1766 ,27322 ,7025 ,10117 ,31213 ,29411 ,23459 ,15623 ,29566 ,
      13949 ,14611 ,5457 ,22703 ,4658 ,1193 ,19750 ,4492 ,25346 ,14545 ,12419 ,23602 ,6308 ,5152 ,4424 ,23295 ,12609 ,8118 ,26599 ,27868 ,25464 ,19967 ,4705 ,21304 ,8723 ,15512 ,9471 ,3766 ,2356 ,17989 ,31325 ,6703 ,13793 ,5773 ,22009 ,12586 ,7559 ,20830 ,26001 ,3275 ,30203 ,17101 ,1240 ,19609 ,29060 ,24393 ,5670 ,24808 ,27265 ,19050 ,20244 ,11031 ,12253 ,19391 ,4532 ,7068 ,23502 ,3315 ,13433 ,31606 ,18599 ,4248 ,8276 ,3482 ,3147 ,31890 ,9868 ,29026 ,20156 ,23050 ,2828 ,30163 ,22372 ,26169 ,30518 ,5161 ,5951 ,22363 ,22469 ,11482 ,31942 ,31826 ,4539 ,13027 ,2410 ,29777 ,10548 ,27792 ,28495 ,23637 ,21795 ,10328 ,22996 ,11145 ,25559 ,4325 ,12203 ,8557 ,18514 ,1664 ,32653 ,4983 ,5365 ,3235 ,7191 ,9953 ,16127 ,15910 ,3599 ,32526 ,19797 ,26678 ,11895 ,20135 ,17364 ,14443 ,16779 ,10624 ,13218 ,18843 ,25858 ,6457 ,24712 ,27979 ,9902 ,10717 ,28432 ,7439 ,12128 ,12952 ,19675 ,19316 ,11916 ,27229 ,15725 ,12379 ,27247 ,30185 ,13931 ,8705 ,31924 ,22354 ,12185 ,25840 ,11934 ,32260 ,27710 ,18676 ,10279 ,15994 ,22094 ,8520 ,6039 ,30654 ,21035 ,28275 ,13164 ,27434 ,5504 ,27304 ,15743 ,2881 ,22750 ,19944 ,8917 ,3774 ,28283 ,1153 ,21433 ,9690 ,7753 ,16043 ,11991 ,13627 ,14877 ,7352 ,12913 ,10062 ,29991 ,24844 ,16953 ,8384 ,23190 ,12041 ,12397 ,2486 ,10408 ,193 ,2239 ,6096 ,2569 ,28626 ,19693 ,9205 ,32156 ,5542 ,30970 ,17535 ,12860 ,25424 ,21247 ,17888 ,15800 ,18433 ,31363 ,22460 ,4918 ,14200 ,7502 ,14345 ,7075 ,17416 ,27516 ,28713 ,28885 ,24186 ,19334 ,32092 ,14658 ,21490 ,3181 ,14044 ,1343 ,29853 ,9811 ,28794 ,32193 ,18131 ,24345 ,29729 ,13996 ,3726 ,12970 ,1543 ,9522 ,3398 ,16206 ,22872 ,30793 ,20401 ,12146 ,6802 ,340 ,26532 ,8823 ,11315 ,28081 ,21621 ,20078 ,12454 ,24036 ,4105 ,730 ,15400 ,20923 ,1033 ,
      18056 ,7427 ,27154 ,23115 ,24733 ,2281 ,26094 ,24637 ,28731 ,9890 ,16995 ,20513 ,23671 ,26669 ,31708 ,22608 ,27534 ,6445 ,25166 ,25582 ,8959 ,6525 ,1366 ,7915 ,6242 ,24700 ,23738 ,12033 ,23921 ,30439 ,22056 ,10963 ,28903 ,14431 ,12633 ,25978 ,20696 ,21669 ,12522 ,31966 ,11958 ,11883 ,697 ,27483 ,6275 ,7526 ,22963 ,16746 ,19570 ,10612 ,14952 ,17137 ,1978 ,30291 ,10321 ,21483 ,24204 ,13206 ,25774 ,16449 ,31098 ,4801 ,20314 ,5230 ,7093 ,3223 ,25144 ,3958 ,1856 ,21329 ,11429 ,27688 ,13332 ,32641 ,18868 ,31036 ,31458 ,3590 ,27558 ,27817 ,31012 ,8545 ,23509 ,14495 ,12066 ,30908 ,25284 ,5889 ,17434 ,18502 ,5820 ,24211 ,28529 ,28129 ,21646 ,31405 ,29148 ,15898 ,9242 ,16248 ,23807 ,17809 ,13840 ,13702 ,14363 ,7179 ,8774 ,4609 ,24387 ,32520 ,13621 ,22866 ,7520 ,32514 ,8865 ,20644 ,9291 ,15093 ,1791 ,29304 ,18930 ,19785 ,24309 ,10811 ,23771 ,772 ,19207 ,10201 ,14676 ,11470 ,16821 ,6375 ,16297 ,13311 ,2699 ,26765 ,16318 ,5939 ,6118 ,6888 ,23954 ,9944 ,25325 ,21226 ,1832 ,26157 ,29329 ,3641 ,410 ,30329 ,7606 ,5914 ,21508 ,30506 ,27085 ,16945 ,32695 ,7940 ,30616 ,13881 ,20198 ,29014 ,4378 ,12563 ,30472 ,2364 ,13172 ,7145 ,32110 ,3135 ,20877 ,9765 ,10362 ,8871 ,15679 ,5993 ,19352 ,23038 ,1407 ,29906 ,32703 ,27047 ,26275 ,23929 ,8096 ,2816 ,6991 ,4028 ,15478 ,26135 ,2452 ,1509 ,8422 ,27780 ,14163 ,29234 ,28000 ,2740 ,25506 ,15017 ,14062 ,2398 ,7647 ,16575 ,447 ,16118 ,23403 ,19429 ,3199 ,31814 ,3322 ,22278 ,26316 ,11363 ,25016 ,6350 ,4700 ,4527 ,10543 ,13213 ,22089 ,23185 ,28880 ,28076 ,1361 ,10316 ,25279 ,1786 ,7601 ,26270 ,25011 ,25052 ,25098 ,28483 ,19161 ,29102 ,25728 ,20650 ,26048 ,6196 ,13394 ,11133 ,30061 ,8638 ,10996 ,18641 ,25057 ,2674 ,29871 ,25547 ,12295 ,18339 ,21829 ,21944 ,7828 ,26927 ,
      15818 ,6691 ,25678 ,11766 ,15200 ,22525 ,3549 ,17253 ,2720 ,2344 ,2261 ,17789 ,11816 ,1655 ,5717 ,12688 ,5796 ,15500 ,12727 ,7259 ,25615 ,2904 ,25103 ,27022 ,18451 ,9459 ,32041 ,10054 ,23030 ,20810 ,27209 ,29709 ,13038 ,27856 ,6577 ,29037 ,808 ,1675 ,14454 ,19853 ,17906 ,12597 ,11042 ,24120 ,27879 ,9297 ,22647 ,22714 ,21265 ,19955 ,24855 ,2956 ,18687 ,6850 ,28488 ,19327 ,17427 ,4693 ,17663 ,5553 ,25199 ,18142 ,26543 ,19468 ,26223 ,4480 ,7893 ,28967 ,6478 ,11836 ,32473 ,8498 ,22478 ,4646 ,24440 ,4433 ,11179 ,12194 ,4927 ,20771 ,31381 ,14599 ,13440 ,18374 ,5033 ,20019 ,19166 ,1484 ,17670 ,5445 ,16876 ,25781 ,3050 ,2180 ,16723 ,13568 ,4936 ,23590 ,17942 ,5726 ,15947 ,9643 ,22825 ,14298 ,27620 ,25334 ,23412 ,32436 ,27567 ,15099 ,30107 ,31717 ,8684 ,5140 ,8332 ,30239 ,26453 ,32346 ,29107 ,6966 ,14218 ,4412 ,20492 ,16554 ,21744 ,24487 ,10492 ,21145 ,18385 ,24796 ,31558 ,28978 ,25879 ,5737 ,30250 ,6632 ,17553 ,29048 ,2967 ,14239 ,7270 ,4974 ,9634 ,11777 ,30988 ,17089 ,3980 ,29186 ,29197 ,11521 ,25733 ,28989 ,11580 ,1228 ,23334 ,29983 ,1399 ,29453 ,12341 ,5297 ,12878 ,12574 ,29917 ,17078 ,3652 ,17997 ,27442 ,6386 ,22289 ,13781 ,28358 ,29245 ,19535 ,1797 ,8649 ,30849 ,14506 ,20818 ,29461 ,3969 ,7948 ,16259 ,20655 ,30447 ,25442 ,25989 ,17148 ,26868 ,25593 ,388 ,20979 ,23126 ,32174 ,7056 ,19656 ,29972 ,21990 ,26580 ,9849 ,17345 ,26786 ,12241 ,20351 ,27353 ,8992 ,5356 ,22816 ,11727 ,30884 ,19038 ,31613 ,11569 ,13517 ,31244 ,26053 ,9740 ,5560 ,20232 ,21875 ,16456 ,29512 ,15299 ,674 ,10148 ,31520 ,31594 ,31539 ,29442 ,6558 ,12708 ,7874 ,8313 ,9223 ,23490 ,27135 ,14933 ,4359 ,29310 ,14144 ,30042 ,19711 ,4236 ,18794 ,12330 ,10889 ,11226 ,6201 ,15654 ,26973 ,8264 ,2625 ,24588 ,22204 ,29597 ,1287 ,3849 ,
      9540 ,28614 ,31653 ,10137 ,23231 ,4153 ,2139 ,18243 ,16842 ,2227 ,2591 ,28324 ,23704 ,18834 ,6957 ,19127 ,13816 ,2474 ,11245 ,29501 ,21001 ,15766 ,13399 ,16093 ,3416 ,10396 ,22135 ,185 ,4020 ,26860 ,7715 ,965 ,12767 ,24832 ,10908 ,20221 ,26702 ,22545 ,28926 ,29646 ,1561 ,12901 ,21558 ,7376 ,13061 ,18936 ,20425 ,24895 ,12988 ,8372 ,12790 ,21864 ,892 ,3097 ,11138 ,14037 ,28122 ,23178 ,2173 ,15292 ,14792 ,16644 ,13480 ,8197 ,13259 ,1141 ,6220 ,11558 ,10738 ,15220 ,23549 ,6017 ,22890 ,8905 ,28195 ,24508 ,30366 ,16770 ,26444 ,5406 ,16224 ,2869 ,18606 ,30873 ,23856 ,14727 ,30066 ,14992 ,25206 ,22738 ,11658 ,31105 ,31741 ,14799 ,10589 ,28678 ,30811 ,16031 ,4746 ,31233 ,29369 ,24919 ,21104 ,26352 ,20582 ,21421 ,18277 ,1447 ,5664 ,19791 ,14871 ,30787 ,22957 ,13615 ,15673 ,26042 ,22641 ,30101 ,8643 ,14138 ,20419 ,14865 ,3362 ,9066 ,4573 ,24084 ,547 ,2053 ,10687 ,25828 ,18813 ,17334 ,9923 ,3569 ,1634 ,5335 ,29747 ,31912 ,4295 ,21765 ,31860 ,20126 ,5131 ,22439 ,24363 ,30173 ,3245 ,21979 ,3285 ,18569 ,11001 ,4502 ,1163 ,13919 ,23265 ,12389 ,8088 ,25434 ,3736 ,31295 ,14014 ,19304 ,24156 ,7045 ,17858 ,31333 ,5512 ,12830 ,11285 ,12116 ,1003 ,24006 ,28764 ,24315 ,3368 ,30763 ,22324 ,27217 ,12349 ,19645 ,30624 ,13134 ,18646 ,22064 ,3744 ,15713 ,7322 ,7723 ,10032 ,16923 ,163 ,2539 ,32211 ,8508 ,14308 ,27342 ,19863 ,17717 ,9418 ,17263 ,6396 ,10267 ,4187 ,6642 ,6741 ,17355 ,8323 ,8459 ,7155 ,32248 ,4255 ,26775 ,20546 ,15027 ,25062 ,22253 ,18149 ,27698 ,13712 ,4808 ,31976 ,16651 ,1955 ,24647 ,12840 ,28263 ,19730 ,5345 ,19243 ,17273 ,17212 ,17202 ,28812 ,6027 ,26362 ,583 ,29656 ,10817 ,9072 ,18253 ,9829 ,27422 ,3529 ,22805 ,11409 ,12502 ,2679 ,24991 ,9398 ,5492 ,2119 ,21084 ,17028 ,3908 ,31183 ,15593 ,
      21914 ,29841 ,2644 ,30031 ,28453 ,25698 ,1756 ,24981 ,11333 ,3169 ,28046 ,10513 ,27750 ,27970 ,16545 ,23373 ,8841 ,32080 ,7115 ,4348 ,2786 ,15448 ,29876 ,26245 ,13281 ,14646 ,21196 ,6088 ,26127 ,380 ,16915 ,30586 ,28099 ,17404 ,5859 ,23479 ,32611 ,31428 ,3928 ,11399 ,15063 ,7490 ,10171 ,24279 ,15868 ,23777 ,4579 ,13591 ,26639 ,28701 ,24607 ,27124 ,24670 ,23891 ,25552 ,1336 ,21639 ,28873 ,16716 ,667 ,10582 ,1948 ,16419 ,20284 ,358 ,25412 ,30417 ,29431 ,13751 ,19505 ,17048 ,27412 ,11491 ,30958 ,5267 ,23304 ,24766 ,25849 ,14209 ,9604 ,29280 ,9193 ,8283 ,31509 ,8234 ,22174 ,12300 ,6171 ,26550 ,32144 ,11697 ,20321 ,19008 ,13487 ,16426 ,644 ,20780 ,18421 ,26992 ,12697 ,2314 ,11786 ,11736 ,3519 ,6820 ,21235 ,19438 ,17633 ,27826 ,778 ,24090 ,22617 ,12164 ,22448 ,8468 ,7863 ,5415 ,3020 ,18344 ,19136 ,9613 ,4906 ,31687 ,23382 ,5110 ,26423 ,16524 ,10462 ,24054 ,20389 ,14108 ,15643 ,21391 ,5634 ,31203 ,21074 ,14697 ,16194 ,28648 ,11628 ,1111 ,10708 ,24478 ,26414 ,18906 ,1531 ,29616 ,10878 ,23148 ,14762 ,21834 ,11108 ,4123 ,9510 ,19097 ,2561 ,2444 ,20971 ,155 ,7685 ,16621 ,18119 ,22223 ,4225 ,10237 ,6711 ,27312 ,9388 ,12472 ,9799 ,15563 ,2089 ,28233 ,19213 ,553 ,9042 ,20096 ,29717 ,5305 ,18783 ,13889 ,8058 ,21949 ,10971 ,31303 ,13984 ,30733 ,973 ,27187 ,30594 ,7693 ,133 ,1918 ,21609 ,1306 ,24577 ,7460 ,15838 ,23449 ,3898 ,15418 ,8811 ,30556 ,21166 ,29811 ,28423 ,10483 ,16515 ,748 ,6790 ,3489 ,26962 ,4876 ,5080 ,7833 ,18314 ,19475 ,328 ,9574 ,5237 ,9163 ,8204 ,20291 ,16396 ,20941 ,4093 ,11078 ,29586 ,16164 ,1081 ,15613 ,31173 ,8028 ,20066 ,103 ,30703 ,18089 ,10207 ,2059 ,523 ,28393 ,15388 ,3868 ,1276 ,298 ,9133 ,26932 ,7803 ,1051 ,20911 ,493 ,73 ,15358 ,268 ,43 ,13 ,
      32765 ,15343 ,20896 ,478 ,1261 ,28378 ,9118 ,26917 ,31158 ,16149 ,4078 ,11063 ,30688 ,8013 ,10192 ,2044 ,16500 ,29796 ,8796 ,30541 ,24562 ,1903 ,15823 ,23434 ,18299 ,4861 ,6775 ,3474 ,5222 ,19460 ,8189 ,20276 ,7670 ,2429 ,9495 ,19082 ,10863 ,18891 ,14747 ,21819 ,21059 ,21376 ,20374 ,14093 ,11613 ,14682 ,10693 ,24463 ,9027 ,28218 ,9784 ,15548 ,4210 ,16606 ,6696 ,27297 ,10956 ,13874 ,29702 ,5290 ,958 ,31288 ,30579 ,7678 ,20269 ,10567 ,28858 ,16701 ,27109 ,26624 ,23876 ,25537 ,11384 ,32596 ,17389 ,5844 ,24264 ,15048 ,23762 ,4564 ,23358 ,27735 ,3154 ,28031 ,30016 ,21899 ,25683 ,1741 ,26230 ,2771 ,32065 ,7100 ,6073 ,13266 ,365 ,16900 ,629 ,18993 ,32129 ,11682 ,31494 ,29265 ,22159 ,12285 ,27397 ,13736 ,25397 ,30402 ,23289 ,11476 ,25834 ,14194 ,22602 ,27811 ,21220 ,19423 ,12682 ,20765 ,11771 ,11721 ,19121 ,5400 ,22433 ,8453 ,23367 ,9598 ,26408 ,16509 ,2038 ,4558 ,14850 ,3347 ,26027 ,22942 ,30086 ,8628 ,26337 ,29354 ,16016 ,4731 ,1432 ,20567 ,19776 ,14856 ,5391 ,30351 ,8890 ,28180 ,11543 ,13244 ,15205 ,23534 ,14977 ,23841 ,2854 ,18591 ,31090 ,25191 ,14784 ,10574 ,950 ,4005 ,10381 ,22120 ,29486 ,13801 ,15751 ,13384 ,18228 ,23216 ,28599 ,31638 ,28309 ,16827 ,18819 ,6942 ,24880 ,13046 ,12886 ,21543 ,20206 ,12752 ,22530 ,28911 ,14022 ,877 ,8357 ,12775 ,15277 ,28107 ,16629 ,13465 ,2524 ,10017 ,15698 ,7307 ,19630 ,22309 ,13119 ,18631 ,12815 ,17843 ,19289 ,24141 ,23991 ,11270 ,24300 ,3353 ,22424 ,31845 ,31897 ,4280 ,17319 ,10672 ,3554 ,1619 ,4487 ,3270 ,30158 ,3230 ,12374 ,1148 ,25419 ,3721 ,24632 ,31961 ,27683 ,13697 ,26760 ,7140 ,15012 ,25047 ,17248 ,19848 ,8493 ,14293 ,6627 ,6381 ,17340 ,8308 ,18238 ,29641 ,6012 ,26347 ,5330 ,12825 ,17258 ,17197 ,24976 ,11394 ,27407 ,3514 ,21069 ,9383 ,3893 ,31168 ,
      26912 ,21814 ,25532 ,12280 ,8623 ,13379 ,18626 ,25042 ,25037 ,7586 ,10301 ,25264 ,29087 ,25083 ,20635 ,26033 ,19414 ,432 ,2383 ,7632 ,29219 ,8407 ,2725 ,25491 ,6335 ,26301 ,31799 ,3307 ,13198 ,4685 ,23170 ,28865 ,13866 ,32680 ,30491 ,27070 ,3626 ,1817 ,30314 ,7591 ,26750 ,16282 ,11455 ,16806 ,6873 ,16303 ,9929 ,25310 ,5978 ,10347 ,3120 ,20862 ,12548 ,20183 ,2349 ,13157 ,23914 ,32688 ,23023 ,1392 ,4013 ,8081 ,26120 ,2437 ,5215 ,31083 ,13191 ,25759 ,17122 ,19555 ,30276 ,10306 ,31951 ,20681 ,14416 ,12618 ,27468 ,11943 ,7511 ,22948 ,22593 ,23656 ,9875 ,16980 ,23100 ,18041 ,2266 ,26079 ,7900 ,8944 ,6430 ,25151 ,12018 ,6227 ,30424 ,22041 ,31390 ,28514 ,18487 ,5805 ,14480 ,30997 ,30893 ,25269 ,27673 ,1841 ,3208 ,25129 ,31021 ,13317 ,3575 ,27543 ,22851 ,24372 ,7164 ,8759 ,16233 ,29133 ,17794 ,13825 ,29289 ,9276 ,32499 ,8850 ,10796 ,18915 ,757 ,19192 ,21130 ,21729 ,4397 ,20477 ,30224 ,8669 ,32331 ,29092 ,14283 ,15932 ,23575 ,17927 ,32421 ,27605 ,15084 ,30092 ,20756 ,11164 ,4631 ,24425 ,28952 ,26208 ,11821 ,32458 ,1469 ,5018 ,14584 ,13425 ,25766 ,17655 ,2165 ,16708 ,29694 ,23015 ,9444 ,32026 ,7244 ,5781 ,2889 ,25088 ,17238 ,15185 ,6676 ,25663 ,17774 ,2705 ,1640 ,5702 ,22699 ,27864 ,12582 ,11027 ,29022 ,13023 ,1660 ,14439 ,19312 ,18672 ,19940 ,24840 ,5538 ,17412 ,18127 ,26528 ,23111 ,25578 ,25974 ,17133 ,3954 ,14491 ,16244 ,20640 ,6371 ,3637 ,12559 ,29902 ,29230 ,22274 ,1782 ,8634 ,11762 ,7255 ,29033 ,2952 ,28963 ,18370 ,5722 ,30235 ,28974 ,29182 ,17074 ,3965 ,29968 ,11565 ,29438 ,12326 ,10133 ,29497 ,20217 ,21860 ,11554 ,30869 ,31229 ,26038 ,17330 ,21975 ,7041 ,19641 ,27338 ,26771 ,5341 ,22801 ,30027 ,4344 ,23475 ,27120 ,29427 ,31505 ,12693 ,7859 ,15639 ,10874 ,4221 ,18779 ,24573 ,26958 ,29582 ,1272 ,
      474 ,30537 ,19078 ,15544 ,16697 ,28027 ,11678 ,19419 ,3343 ,28176 ,22116 ,21539 ,7303 ,4276 ,13693 ,26343 ,12276 ,7628 ,27066 ,20858 ,25755 ,16976 ,5801 ,8755 ,20473 ,24421 ,32022 ,11023 ,17129 ,2948 ,21856 ,27116 ,15540 ,20854 ,32722 ,32726 ,5007 ,18017 ,2001 ,437 ,23981 ,7971 ,8146 ,3798 ,18710 ,16324 ,29753 ,19995 ,10098 ,5180 ,915 ,32730 ,14573 ,28576 ,15505 ,30647 ,24693 ,30499 ,9452 ,1221 ,10389 ,13912 ,14639 ,9503 ,4854 ,23834 ,26294 ,5011 ,24414 ,3672 ,8585 ,2388 ,17833 ,32554 ,15162 ,9318 ,9981 ,21693 ,23798 ,29360 ,31485 ,26188 ,20163 ,18021 ,20745 ,1883 ,12732 ,10652 ,6485 ,1699 ,28556 ,1863 ,9667 ,10745 ,13758 ,12093 ,24943 ,22391 ,18195 ,2005 ,26197 ,22569 ,31125 ,7637 ,19279 ,20723 ,17297 ,23078 ,6302 ,5945 ,31918 ,31357 ,23665 ,31452 ,23948 ,441 ,11810 ,11173 ,7264 ,8986 ,23698 ,30360 ,31854 ,6735 ,27744 ,24760 ,1105 ,29805 ,30682 ,24258 ,1426 ,23985 ,29081 ,27462 ,32415 ,29224 ,7297 ,9975 ,32288 ,27900 ,32294 ,25906 ,15889 ,16022 ,18984 ,22382 ,7201 ,7975 ,30213 ,1719 ,25620 ,25356 ,21443 ,3679 ,19897 ,27257 ,19562 ,21257 ,12980 ,26631 ,9019 ,5970 ,10090 ,8150 ,21718 ,22017 ,22758 ,8412 ,2514 ,9341 ,29539 ,16349 ,17586 ,6124 ,4301 ,13544 ,26821 ,6585 ,29925 ,3802 ,4386 ,6919 ,2909 ,12641 ,24164 ,13655 ,25931 ,10916 ,9718 ,5867 ,22231 ,6149 ,5597 ,22488 ,27630 ,18714 ,17916 ,17481 ,25226 ,2730 ,22299 ,835 ,17751 ,17563 ,27906 ,26796 ,9233 ,4737 ,32120 ,18186 ,23057 ,16328 ,14272 ,14072 ,25108 ,25642 ,11843 ,13342 ,14373 ,21336 ,11968 ,15227 ,19512 ,28741 ,11295 ,15974 ,19371 ,29757 ,27594 ,6406 ,28822 ,25496 ,13109 ,22900 ,20592 ,26480 ,1571 ,6894 ,21771 ,16852 ,11206 ,11501 ,6830 ,19999 ,15073 ,6505 ,27027 ,11343 ,12482 ,18549 ,3077 ,14707 ,3000 ,15428 ,8038 ,5060 ,
      29551 ,29396 ,7010 ,10102 ,5691 ,29937 ,25943 ,6340 ,1609 ,7213 ,19909 ,22668 ,32300 ,32390 ,4600 ,1438 ,30393 ,23069 ,14385 ,5184 ,17763 ,10765 ,18456 ,27642 ,20604 ,8592 ,31768 ,19383 ,30283 ,6842 ,3089 ,23883 ,16598 ,20175 ,28568 ,919 ,15174 ,31059 ,14819 ,26306 ,17309 ,26729 ,27376 ,18207 ,13088 ,23960 ,31866 ,4456 ,8158 ,24531 ,4047 ,32734 ,6665 ,927 ,9464 ,21028 ,23731 ,27078 ,32034 ,23327 ,22128 ,23258 ,21189 ,19090 ,6768 ,2847 ,31792 ,14577 ,32015 ,19890 ,31761 ,31804 ,31835 ,15143 ,32003 ,8127 ,25912 ,32269 ,14354 ,20573 ,27388 ,19270 ,2835 ,28580 ,29683 ,4059 ,32046 ,25378 ,32480 ,14397 ,31780 ,11436 ,19921 ,23556 ,17055 ,7022 ,14608 ,14542 ,8115 ,15509 ,5770 ,17098 ,19047 ,3312 ,31887 ,26166 ,31823 ,23634 ,8554 ,9950 ,20132 ,6454 ,12949 ,30182 ,32257 ,30651 ,2878 ,9687 ,10059 ,2483 ,9202 ,17885 ,14342 ,32089 ,28791 ,1540 ,6799 ,12451 ,7424 ,9887 ,6442 ,24697 ,14428 ,11880 ,10609 ,13203 ,3220 ,32638 ,8542 ,18499 ,15895 ,7176 ,32511 ,19782 ,11467 ,5936 ,26154 ,30503 ,29011 ,3132 ,23035 ,2813 ,27777 ,2395 ,31811 ,4524 ,10313 ,28480 ,11130 ,25544 ,6688 ,2341 ,15497 ,9456 ,27853 ,12594 ,19952 ,4690 ,4477 ,4643 ,14596 ,5442 ,23587 ,25331 ,5137 ,4409 ,24793 ,29045 ,17086 ,1225 ,12571 ,13778 ,20815 ,25986 ,7053 ,12238 ,19035 ,20229 ,31591 ,23487 ,4233 ,8261 ,28611 ,2224 ,2471 ,10393 ,24829 ,12898 ,8369 ,23175 ,1138 ,8902 ,2866 ,22735 ,16028 ,21418 ,13612 ,14862 ,25825 ,31909 ,30170 ,13916 ,19301 ,12113 ,27214 ,15710 ,8505 ,10264 ,32245 ,27695 ,28260 ,6024 ,27419 ,5489 ,29838 ,3166 ,32077 ,14643 ,17401 ,7487 ,28698 ,28870 ,25409 ,30955 ,9190 ,32141 ,18418 ,21232 ,22445 ,4903 ,20386 ,16191 ,1528 ,9507 ,18116 ,9796 ,29714 ,13981 ,21606 ,8808 ,6787 ,325 ,4090 ,20063 ,15385 ,20908 ,
      15340 ,16146 ,29793 ,4858 ,2426 ,21373 ,28215 ,13871 ,10564 ,32593 ,27732 ,2768 ,18990 ,13733 ,27808 ,5397 ,4555 ,29351 ,30348 ,23838 ,4002 ,23213 ,13043 ,874 ,10014 ,17840 ,31842 ,3267 ,31958 ,19845 ,29638 ,11391 ,21811 ,7583 ,429 ,26298 ,32677 ,16279 ,10344 ,32685 ,31080 ,20678 ,23653 ,8941 ,28511 ,1838 ,24369 ,9273 ,21726 ,15929 ,11161 ,5015 ,23012 ,15182 ,27861 ,18669 ,25575 ,3634 ,7252 ,29179 ,29494 ,21972 ,4341 ,10871 ,30534 ,28173 ,7625 ,24418 ,20851 ,7968 ,5177 ,30496 ,23831 ,32551 ,26185 ,1696 ,22388 ,20720 ,31449 ,30357 ,24255 ,9972 ,22379 ,3676 ,5967 ,9338 ,6582 ,13652 ,22485 ,832 ,18183 ,13339 ,15971 ,22897 ,11498 ,18546 ,29393 ,7210 ,23066 ,8589 ,20172 ,26726 ,24528 ,27075 ,2844 ,15140 ,19267 ,14394 ,14539 ,26163 ,30179 ,17882 ,9884 ,32635 ,5933 ,2392 ,2338 ,4640 ,29042 ,12235 ,2221 ,8899 ,31906 ,10261 ,3163 ,30952 ,16188 ,8805 ,16143 ,32590 ,29348 ,17837 ,7580 ,20675 ,15926 ,3631 ,28170 ,32548 ,9969 ,829 ,7207 ,15137 ,32632 ,8896 ,32587 ,32545 ,32542 ,32558 ,3615 ,32574 ,813 ,15121 ,19813 ,32561 ,15150 ,7551 ,20688 ,800 ,26694 ,32603 ,10855 ,3618 ,4999 ,15166 ,32669 ,7567 ,8925 ,1822 ,5381 ,32577 ,4842 ,21357 ,858 ,29335 ,3251 ,19829 ,18530 ,816 ,3660 ,9322 ,30480 ,28157 ,1680 ,20704 ,17866 ,15124 ,8573 ,26710 ,12219 ,32619 ,10245 ,30936 ,9351 ,19816 ,10640 ,9985 ,16795 ,845 ,22910 ,30319 ,13234 ,32564 ,20733 ,18961 ,7981 ,4829 ,18859 ,28186 ,17380 ,15153 ,26176 ,21697 ,26739 ,10842 ,14459 ,7223 ,4653 ,7554 ,20151 ,32648 ,11911 ,8912 ,30965 ,24340 ,24728 ,20691 ,1851 ,23802 ,16292 ,30467 ,27995 ,7596 ,15195 ,803 ,6473 ,15942 ,25874 ,3647 ,21985 ,6553 ,23226 ,26697 ,10733 ,29364 ,9918 ,17853 ,19858 ,19238 ,28448 ,32606 ,13746 ,2309 ,21386 ,10232 ,7455 ,16159 ,
      1256 ,10858 ,27104 ,31489 ,26022 ,29481 ,19625 ,26755 ,8618 ,3621 ,17117 ,14475 ,30219 ,7239 ,3949 ,11549 ,16692 ,5002 ,24409 ,26192 ,29076 ,21713 ,17911 ,27589 ,5686 ,15169 ,32010 ,5765 ,14423 ,27848 ,24824 ,17396 ,2421 ,32672 ,20846 ,20167 ,7575 ,32664 ,16790 ,16287 ,26017 ,7570 ,12264 ,13363 ,25475 ,416 ,3291 ,4669 ,22025 ,8928 ,16964 ,18025 ,10290 ,31067 ,12602 ,11927 ,27527 ,1825 ,5789 ,30981 ,13809 ,24356 ,8834 ,18899 ,16493 ,5384 ,19407 ,20749 ,12269 ,18977 ,30386 ,11460 ,4548 ,32580 ,16685 ,26608 ,1725 ,27719 ,7084 ,13250 ,20260 ,4845 ,30525 ,1887 ,26901 ,15327 ,11047 ,7997 ,24447 ,21360 ,19066 ,18875 ,27281 ,28202 ,5274 ,31272 ,13449 ,861 ,21527 ,12736 ,13368 ,3989 ,31622 ,16811 ,14840 ,29338 ,3331 ,22926 ,23518 ,30335 ,18575 ,25175 ,3705 ,3254 ,4264 ,10656 ,18615 ,10001 ,24125 ,11254 ,8292 ,19832 ,13681 ,7124 ,17181 ,29625 ,3498 ,9367 ,5044 ,18533 ,19983 ,6489 ,25480 ,15958 ,26464 ,6878 ,4721 ,819 ,18698 ,17465 ,25626 ,18170 ,21320 ,15211 ,26615 ,3663 ,7959 ,1703 ,29208 ,24242 ,27884 ,25890 ,13528 ,9325 ,8134 ,22001 ,12625 ,6569 ,10900 ,5851 ,9487 ,30483 ,32714 ,28560 ,421 ,20838 ,3782 ,16308 ,26327 ,28160 ,15528 ,28011 ,8739 ,7612 ,11007 ,2932 ,12077 ,1683 ,18005 ,1867 ,2372 ,23818 ,9302 ,21677 ,31341 ,20707 ,1989 ,22553 ,8970 ,31436 ,6719 ,24744 ,12435 ,17869 ,30635 ,9671 ,3296 ,14526 ,23618 ,9934 ,20557 ,15127 ,14561 ,19874 ,25362 ,19254 ,11420 ,23540 ,23867 ,8576 ,5168 ,10749 ,6324 ,29380 ,22652 ,32374 ,4440 ,26713 ,903 ,31043 ,21012 ,24515 ,23311 ,23242 ,8245 ,12222 ,1209 ,13762 ,4674 ,2325 ,5426 ,25315 ,19766 ,32622 ,24681 ,11864 ,2797 ,5920 ,4508 ,28464 ,5473 ,10248 ,13900 ,12097 ,23159 ,2208 ,22719 ,21402 ,4887 ,30939 ,14627 ,7471 ,13965 ,16175 ,309 ,20047 ,
      7769 ,9354 ,6137 ,24947 ,22030 ,17168 ,16059 ,5983 ,6932 ,19819 ,9706 ,6598 ,21449 ,13668 ,5880 ,14983 ,1732 ,10643 ,13643 ,22395 ,12007 ,3692 ,21270 ,30129 ,14893 ,9988 ,25919 ,19601 ,27475 ,24112 ,7368 ,24271 ,14085 ,16798 ,3790 ,18199 ,8933 ,13355 ,15240 ,10352 ,28299 ,848 ,26809 ,15248 ,17494 ,21514 ,1169 ,22501 ,22766 ,22913 ,6907 ,2009 ,6419 ,14827 ,19960 ,15987 ,6518 ,30322 ,2897 ,11514 ,15759 ,18562 ,15441 ,14755 ,1896 ,13237 ,8400 ,26201 ,16969 ,1712 ,10758 ,3125 ,23206 ,32567 ,21706 ,24235 ,3685 ,16672 ,12057 ,23847 ,30007 ,20736 ,5958 ,22573 ,22582 ,16480 ,24860 ,22404 ,11186 ,18964 ,10078 ,31465 ,12929 ,30373 ,24773 ,25805 ,10424 ,7984 ,16337 ,31129 ,18030 ,26888 ,209 ,20867 ,28589 ,4832 ,2502 ,5193 ,12413 ,30512 ,13925 ,15794 ,16989 ,18862 ,6112 ,7641 ,2255 ,24434 ,2961 ,20345 ,2585 ,28189 ,4289 ,4181 ,28040 ,5261 ,28642 ,30550 ,4072 ,17383 ,16010 ,19283 ,10295 ,14410 ,23569 ,12553 ,22110 ,15156 ,32282 ,17745 ,19903 ,31997 ,8536 ,2860 ,27726 ,26179 ,9963 ,20727 ,17111 ,16679 ,18692 ,14555 ,9700 ,21700 ,32276 ,30195 ,11950 ,17898 ,1553 ,15055 ,21051 ,26742 ,23973 ,17301 ,31072 ,26009 ,28291 ,20188 ,940 ,10845 ,30670 ,24544 ,6055 ,27091 ,23271 ,12664 ,10778 ,14462 ,27450 ,23082 ,13180 ,8605 ,6855 ,12530 ,5520 ,7226 ,32403 ,28934 ,29950 ,3936 ,27320 ,29409 ,13947 ,4656 ,25344 ,6306 ,12607 ,25462 ,8721 ,2354 ,13791 ,7557 ,30201 ,29058 ,27263 ,12251 ,23500 ,18597 ,3145 ,20154 ,22370 ,5949 ,31940 ,2408 ,28493 ,22994 ,12201 ,32651 ,7189 ,3597 ,11893 ,16777 ,25856 ,9900 ,12126 ,11914 ,27245 ,31922 ,11932 ,10277 ,6037 ,13162 ,15741 ,8915 ,21431 ,11989 ,12911 ,16951 ,12395 ,2237 ,19691 ,30968 ,21245 ,31361 ,7500 ,27514 ,19332 ,3179 ,9809 ,24343 ,12968 ,16204 ,12144 ,8821 ,20076 ,728 ,
      18054 ,24731 ,28729 ,23669 ,27532 ,8957 ,6240 ,23919 ,28901 ,20694 ,11956 ,6273 ,19568 ,1976 ,24202 ,31096 ,7091 ,1854 ,13330 ,31456 ,31010 ,12064 ,17432 ,28527 ,29146 ,23805 ,14361 ,24385 ,7518 ,9289 ,18928 ,23769 ,14674 ,16295 ,16316 ,23952 ,1830 ,408 ,21506 ,32693 ,20196 ,30470 ,32108 ,10360 ,19350 ,32701 ,8094 ,15476 ,8420 ,27998 ,14060 ,445 ,3197 ,26314 ,4698 ,22087 ,1359 ,7599 ,25096 ,25726 ,13392 ,10994 ,29869 ,21827 ,15816 ,15198 ,2718 ,11814 ,5794 ,25613 ,18449 ,23028 ,13036 ,806 ,17904 ,27877 ,21263 ,18685 ,17425 ,25197 ,26221 ,6476 ,22476 ,11177 ,31379 ,5031 ,17668 ,3048 ,4934 ,15945 ,27618 ,27565 ,8682 ,26451 ,14216 ,21742 ,18383 ,25877 ,17551 ,7268 ,30986 ,29195 ,11578 ,1397 ,12876 ,3650 ,22287 ,19533 ,14504 ,7946 ,25440 ,25591 ,32172 ,21988 ,26784 ,8990 ,30882 ,13515 ,5558 ,29510 ,31518 ,6556 ,9221 ,4357 ,19709 ,10887 ,26971 ,22202 ,9538 ,23229 ,16840 ,23702 ,13814 ,20999 ,3414 ,4018 ,12765 ,26700 ,1559 ,13059 ,12986 ,890 ,28120 ,14790 ,13257 ,10736 ,22888 ,30364 ,16222 ,23854 ,25204 ,31739 ,30809 ,29367 ,20580 ,5662 ,22955 ,22639 ,20417 ,4571 ,10685 ,9921 ,29745 ,31858 ,24361 ,3283 ,1161 ,8086 ,14012 ,17856 ,11283 ,28762 ,22322 ,30622 ,3742 ,10030 ,32209 ,19861 ,6394 ,6739 ,7153 ,20544 ,18147 ,31974 ,12838 ,19241 ,28810 ,29654 ,9827 ,11407 ,9396 ,17026 ,21912 ,28451 ,11331 ,27748 ,8839 ,2784 ,13279 ,26125 ,28097 ,32609 ,15061 ,15866 ,26637 ,24668 ,21637 ,10580 ,356 ,13749 ,11489 ,24764 ,29278 ,8232 ,26548 ,19006 ,20778 ,2312 ,6818 ,27824 ,12162 ,5413 ,9611 ,5108 ,24052 ,21389 ,14695 ,1109 ,18904 ,23146 ,4121 ,2442 ,16619 ,10235 ,12470 ,28231 ,20094 ,13887 ,31301 ,27185 ,1916 ,7458 ,15416 ,29809 ,746 ,4874 ,19473 ,9161 ,20939 ,16162 ,8026 ,18087 ,28391 ,296 ,1049 ,15356 ,
      32763 ,1259 ,31156 ,30686 ,16498 ,24560 ,18297 ,5220 ,7668 ,10861 ,21057 ,11611 ,9025 ,4208 ,10954 ,956 ,20267 ,27107 ,11382 ,24262 ,23356 ,30014 ,26228 ,6071 ,627 ,31492 ,27395 ,23287 ,22600 ,12680 ,19119 ,23365 ,2036 ,26025 ,26335 ,1430 ,5389 ,11541 ,14975 ,31088 ,948 ,29484 ,18226 ,28307 ,24878 ,20204 ,14020 ,15275 ,2522 ,19628 ,12813 ,23989 ,22422 ,17317 ,4485 ,12372 ,24630 ,26758 ,17246 ,6625 ,18236 ,5328 ,24974 ,21067 ,26910 ,8621 ,25035 ,29085 ,19412 ,29217 ,6333 ,13196 ,13864 ,3624 ,26748 ,6871 ,5976 ,12546 ,23912 ,4011 ,5213 ,17120 ,31949 ,27466 ,22591 ,23098 ,7898 ,12016 ,31388 ,14478 ,27671 ,31019 ,22849 ,16231 ,29287 ,10794 ,21128 ,30222 ,14281 ,32419 ,20754 ,28950 ,1467 ,25764 ,29692 ,7242 ,17236 ,17772 ,22697 ,29020 ,19310 ,5536 ,23109 ,3952 ,6369 ,29228 ,11760 ,28961 ,28972 ,29966 ,10131 ,11552 ,17328 ,27336 ,30025 ,29425 ,15637 ,24571 ,472 ,16695 ,3341 ,7301 ,12274 ,25753 ,20471 ,17127 ,15538 ,5005 ,23979 ,18708 ,10096 ,14571 ,24691 ,10387 ,4852 ,24412 ,17831 ,9979 ,31483 ,20743 ,6483 ,9665 ,24941 ,26195 ,19277 ,6300 ,23663 ,11808 ,23696 ,27742 ,30680 ,29079 ,7295 ,32292 ,18982 ,30211 ,21441 ,19560 ,9017 ,21716 ,2512 ,17584 ,26819 ,4384 ,24162 ,9716 ,5595 ,17914 ,22297 ,27904 ,32118 ,14270 ,11841 ,11966 ,11293 ,27592 ,13107 ,1569 ,11204 ,15071 ,12480 ,2998 ,29549 ,5689 ,1607 ,32298 ,30391 ,17761 ,20602 ,30281 ,16596 ,15172 ,17307 ,13086 ,8156 ,6663 ,23729 ,22126 ,6766 ,32013 ,31833 ,25910 ,27386 ,29681 ,32478 ,19919 ,14606 ,5768 ,31885 ,8552 ,12947 ,2876 ,9200 ,28789 ,7422 ,14426 ,3218 ,15893 ,11465 ,29009 ,27775 ,10311 ,6686 ,27851 ,4475 ,23585 ,24791 ,12569 ,7051 ,31589 ,28609 ,24827 ,1136 ,16026 ,25823 ,19299 ,8503 ,28258 ,29836 ,17399 ,25407 ,18416 ,20384 ,18114 ,21604 ,4088 ,
      15338 ,2424 ,10562 ,18988 ,4553 ,4000 ,10012 ,31956 ,21809 ,32675 ,31078 ,28509 ,21724 ,23010 ,25573 ,29492 ,30532 ,20849 ,23829 ,22386 ,24253 ,5965 ,22483 ,15969 ,29391 ,20170 ,2842 ,14537 ,9882 ,2336 ,2219 ,3161 ,16141 ,7578 ,28168 ,7205 ,32585 ,3613 ,19811 ,20686 ,10853 ,32667 ,5379 ,856 ,18528 ,30478 ,17864 ,12217 ,9349 ,16793 ,13232 ,7979 ,17378 ,26737 ,4651 ,11909 ,24726 ,16290 ,15193 ,25872 ,23224 ,9916 ,28446 ,21384 ,1254 ,26020 ,8616 ,30217 ,16690 ,29074 ,5684 ,14421 ,2419 ,7573 ,26015 ,25473 ,22023 ,10288 ,27525 ,13807 ,16491 ,12267 ,4546 ,1723 ,20258 ,26899 ,24445 ,27279 ,13447 ,13366 ,14838 ,23516 ,3703 ,18613 ,8290 ,17179 ,5042 ,25478 ,4719 ,25624 ,26613 ,29206 ,13526 ,12623 ,9485 ,419 ,26325 ,8737 ,12075 ,2370 ,31339 ,8968 ,12433 ,3294 ,20555 ,25360 ,23865 ,6322 ,4438 ,21010 ,8243 ,4672 ,19764 ,2795 ,5471 ,23157 ,4885 ,13963 ,7767 ,22028 ,6930 ,21447 ,1730 ,12005 ,14891 ,27473 ,14083 ,8931 ,28297 ,17492 ,22764 ,6417 ,6516 ,15757 ,1894 ,16967 ,23204 ,3683 ,30005 ,22580 ,11184 ,12927 ,10422 ,18028 ,28587 ,12411 ,16987 ,2253 ,2583 ,28038 ,4070 ,10293 ,22108 ,19901 ,27724 ,17109 ,9698 ,11948 ,21049 ,31070 ,938 ,6053 ,10776 ,13178 ,5518 ,29948 ,13945 ,12605 ,13789 ,27261 ,3143 ,31938 ,12199 ,11891 ,12124 ,11930 ,15739 ,12909 ,19689 ,7498 ,9807 ,12142 ,18052 ,27530 ,28899 ,19566 ,7089 ,31008 ,29144 ,7516 ,14672 ,1828 ,20194 ,19348 ,8418 ,3195 ,1357 ,13390 ,15814 ,5792 ,13034 ,21261 ,26219 ,31377 ,4932 ,8680 ,18381 ,30984 ,12874 ,14502 ,32170 ,30880 ,31516 ,19707 ,9536 ,13812 ,12763 ,12984 ,13255 ,16220 ,30807 ,22953 ,10683 ,24359 ,14010 ,22320 ,32207 ,7151 ,12836 ,9825 ,21910 ,8837 ,28095 ,26635 ,354 ,29276 ,20776 ,12160 ,24050 ,18902 ,16617 ,20092 ,1914 ,744 ,20937 ,28389 ,
      32761 ,16496 ,7666 ,9023 ,20265 ,23354 ,625 ,22598 ,2034 ,5387 ,946 ,24876 ,2520 ,22420 ,24628 ,18234 ,26908 ,19410 ,13862 ,5974 ,5211 ,22589 ,31386 ,22847 ,21126 ,20752 ,29690 ,22695 ,23107 ,11758 ,10129 ,30023 ,470 ,12272 ,15536 ,10094 ,4850 ,31481 ,24939 ,23661 ,30678 ,18980 ,9015 ,26817 ,5593 ,32116 ,11291 ,11202 ,29547 ,30389 ,16594 ,8154 ,6764 ,27384 ,14604 ,12945 ,7420 ,11463 ,6684 ,24789 ,28607 ,25821 ,29834 ,20382 ,15336 ,4551 ,21807 ,21722 ,30530 ,24251 ,29389 ,9880 ,16139 ,32583 ,10851 ,18526 ,9347 ,17376 ,24724 ,23222 ,1252 ,16688 ,2417 ,22021 ,16489 ,20256 ,13445 ,3701 ,5040 ,26611 ,9483 ,12073 ,12431 ,23863 ,8241 ,5469 ,7765 ,1728 ,14081 ,22762 ,1892 ,30003 ,10420 ,16985 ,4068 ,27722 ,21047 ,10774 ,13943 ,3141 ,12122 ,19687 ,18050 ,7087 ,14670 ,8416 ,15812 ,26217 ,18379 ,32168 ,9534 ,13253 ,10681 ,32205 ,21908 ,352 ,24048 ,1912 ,32759 ,20263 ,2032 ,2518 ,26906 ,5209 ,21124 ,23105 ,468 ,4848 ,30676 ,5591 ,29545 ,6762 ,7418 ,28605 ,15334 ,30528 ,16137 ,9345 ,1250 ,16487 ,5038 ,12429 ,7763 ,1890 ,4066 ,13941 ,18048 ,15810 ,9532 ,21906 ,32757 ,26904 ,466 ,29543 ,15332 ,1248 ,7761 ,18046 ,32755 ,15330 ,32753 ,225 ,227 ,20883 ,1009 ,3825 ,229 ,11050 ,28366 ,16353 ,20885 ,31145 ,20024 ,705 ,1011 ,8000 ,9106 ,21566 ,3827 ,10179 ,15571 ,10440 ,231 ,24450 ,23422 ,17590 ,11052 ,11600 ,18741 ,2271 ,28368 ,21363 ,24550 ,2977 ,16355 ,20361 ,27145 ,31644 ,20887 ,19069 ,29784 ,6128 ,31147 ,7657 ,19171 ,26507 ,20026 ,18878 ,8784 ,30915 ,707 ,14734 ,22181 ,17005 ,1013 ,27284 ,3462 ,4305 ,8002 ,4197 ,26372 ,26084 ,9108 ,28205 ,18287 ,27927 ,21568 ,9771 ,24012 ,2601 ,3829 ,5277 ,19448 ,13548 ,10181 ,10943 ,1489 ,28056 ,15573 ,31275 ,8177 ,28658 ,10442 ,30566 ,113 ,16376 ,
      233 ,13452 ,16888 ,26825 ,24452 ,15264 ,4766 ,7905 ,23424 ,864 ,6061 ,17954 ,17592 ,8344 ,20504 ,28315 ,11054 ,21530 ,2759 ,6589 ,11602 ,24867 ,17675 ,17510 ,18743 ,12739 ,32053 ,1185 ,2273 ,22517 ,4145 ,25690 ,28370 ,13371 ,28019 ,29929 ,21365 ,29473 ,17160 ,8949 ,24552 ,3992 ,23346 ,15256 ,2979 ,10368 ,28770 ,31570 ,16357 ,31625 ,21887 ,3806 ,20363 ,18215 ,5450 ,19668 ,27147 ,16814 ,25671 ,31551 ,31646 ,18806 ,2637 ,14101 ,20889 ,14843 ,25525 ,4390 ,19071 ,1419 ,7003 ,6435 ,29786 ,29341 ,27097 ,19976 ,6130 ,16003 ,28722 ,16833 ,31149 ,3334 ,10555 ,6923 ,7659 ,2025 ,16881 ,14175 ,19173 ,22929 ,28846 ,25291 ,26509 ,30073 ,12307 ,22782 ,20028 ,23521 ,5832 ,2913 ,18880 ,11530 ,31253 ,25156 ,8786 ,30338 ,11372 ,9254 ,30917 ,8877 ,24321 ,6534 ,709 ,18578 ,15036 ,12645 ,14736 ,14964 ,25786 ,15775 ,22183 ,25178 ,23750 ,15457 ,17007 ,14771 ,5089 ,27166 ,1015 ,3708 ,14182 ,24168 ,27286 ,12361 ,7334 ,12023 ,3464 ,3257 ,23277 ,21286 ,4307 ,30145 ,26660 ,18825 ,8004 ,4267 ,13724 ,13659 ,4199 ,22411 ,3055 ,14320 ,26374 ,10659 ,25385 ,19742 ,26086 ,3541 ,2131 ,1748 ,9110 ,18618 ,11670 ,25935 ,28207 ,19617 ,16051 ,6232 ,18289 ,10004 ,617 ,4758 ,27929 ,15685 ,3374 ,14909 ,21570 ,24128 ,29253 ,10920 ,9773 ,12802 ,2185 ,27491 ,24014 ,11257 ,22147 ,7384 ,2603 ,24287 ,2097 ,31665 ,3831 ,8295 ,11709 ,9722 ,5279 ,6614 ,30831 ,30429 ,19450 ,19835 ,12670 ,27004 ,13550 ,8480 ,31699 ,6948 ,10183 ,13684 ,27799 ,5871 ,10945 ,24619 ,16728 ,21465 ,1491 ,7127 ,21208 ,5896 ,28058 ,14999 ,6178 ,2656 ,15575 ,17184 ,8441 ,22235 ,31277 ,5317 ,30745 ,22046 ,8179 ,29628 ,19109 ,16075 ,28660 ,5999 ,30769 ,14120 ,10444 ,3501 ,9586 ,6153 ,30568 ,24963 ,13573 ,1318 ,115 ,9370 ,26396 ,11090 ,16378 ,3880 ,505 ,7785 ,
      235 ,5047 ,19180 ,5601 ,13454 ,2987 ,27937 ,31395 ,16890 ,18536 ,10784 ,17684 ,26827 ,3064 ,16737 ,24886 ,24454 ,19986 ,9264 ,22492 ,15266 ,11193 ,4941 ,17964 ,4768 ,6492 ,32487 ,21296 ,7907 ,27014 ,16085 ,26237 ,23426 ,25483 ,8747 ,27634 ,866 ,27581 ,30121 ,28519 ,6063 ,15961 ,22839 ,17502 ,17956 ,19358 ,22330 ,4950 ,17594 ,26467 ,29121 ,18718 ,8346 ,13096 ,23595 ,8698 ,20506 ,6881 ,17782 ,14232 ,28317 ,21758 ,10506 ,11621 ,11056 ,4724 ,25257 ,17920 ,21532 ,27893 ,22661 ,18492 ,2761 ,822 ,14468 ,17458 ,6591 ,17738 ,6266 ,13052 ,11604 ,18701 ,28502 ,17485 ,24869 ,5584 ,17947 ,21279 ,17677 ,17468 ,18475 ,17441 ,17512 ,25213 ,26557 ,17694 ,18745 ,25629 ,25117 ,25230 ,12741 ,14259 ,3440 ,5810 ,32055 ,18173 ,27661 ,18465 ,1187 ,23044 ,27223 ,17529 ,2275 ,21323 ,13305 ,2734 ,22519 ,11830 ,5731 ,26574 ,4147 ,15214 ,3563 ,17711 ,25692 ,19499 ,5628 ,15832 ,28372 ,26618 ,22936 ,22303 ,13373 ,19549 ,8663 ,14485 ,28021 ,3666 ,27456 ,17475 ,29931 ,19884 ,11874 ,12892 ,21367 ,7962 ,20669 ,839 ,29475 ,18971 ,15952 ,14520 ,17162 ,1706 ,14404 ,25456 ,8951 ,25607 ,20993 ,2778 ,24554 ,29211 ,25747 ,17755 ,3994 ,29068 ,11999 ,31002 ,23348 ,24245 ,5203 ,11594 ,15258 ,1413 ,12355 ,6608 ,2981 ,27887 ,19543 ,17567 ,10370 ,7284 ,9648 ,6283 ,28772 ,25893 ,30264 ,13069 ,31572 ,15876 ,28241 ,18399 ,16359 ,13531 ,26067 ,27910 ,31627 ,17573 ,26490 ,30898 ,21889 ,9328 ,23088 ,5574 ,3808 ,29526 ,688 ,21549 ,20365 ,8137 ,23644 ,26800 ,18217 ,9006 ,22830 ,22678 ,5452 ,22004 ,9863 ,18509 ,19670 ,22745 ,32151 ,32188 ,27149 ,12628 ,25139 ,9237 ,16816 ,4373 ,14158 ,25274 ,25673 ,6572 ,7888 ,17937 ,31553 ,29912 ,19651 ,31534 ,31648 ,10903 ,6215 ,4741 ,18808 ,24151 ,14303 ,19725 ,2639 ,5854 ,30412 ,26987 ,14103 ,22218 ,1301 ,11073 ,
      20891 ,9490 ,28853 ,32124 ,14845 ,10376 ,15693 ,27678 ,25527 ,30486 ,13186 ,18482 ,4392 ,9439 ,25969 ,20212 ,19073 ,32717 ,26289 ,18190 ,1421 ,10085 ,27625 ,19366 ,7005 ,28563 ,31787 ,8110 ,6437 ,15492 ,2466 ,32072 ,29788 ,424 ,7620 ,23061 ,29343 ,4994 ,10635 ,1846 ,27099 ,20841 ,19402 ,21522 ,19978 ,32709 ,30630 ,1204 ,6132 ,3785 ,8395 ,16332 ,16005 ,23968 ,25339 ,27240 ,28724 ,16311 ,2713 ,17546 ,16835 ,29740 ,11326 ,14690 ,31151 ,26330 ,25030 ,14276 ,3336 ,7290 ,1602 ,3213 ,10557 ,28163 ,8611 ,4714 ,6925 ,22103 ,28894 ,12758 ,7661 ,15531 ,21802 ,14076 ,2027 ,461 ,23417 ,3457 ,16883 ,28014 ,25520 ,5827 ,14177 ,11665 ,11704 ,8436 ,19175 ,8742 ,25252 ,25112 ,22931 ,25742 ,26062 ,25134 ,28848 ,7615 ,25025 ,25247 ,25293 ,27053 ,13140 ,1375 ,26511 ,11010 ,25071 ,25646 ,30075 ,20460 ,32441 ,13408 ,12309 ,2935 ,20623 ,29885 ,22784 ,21843 ,7842 ,18762 ,20030 ,12080 ,25298 ,11847 ,23523 ,9654 ,32357 ,31026 ,5834 ,1686 ,6861 ,17448 ,2915 ,28543 ,21660 ,22536 ,18882 ,18008 ,16270 ,13346 ,11532 ,31472 ,27572 ,5748 ,31255 ,1870 ,11443 ,26591 ,25158 ,12719 ,11237 ,7107 ,8788 ,2375 ,27058 ,14377 ,30340 ,24401 ,13635 ,13322 ,11374 ,23821 ,13854 ,2751 ,9256 ,26281 ,18652 ,29162 ,30919 ,9305 ,1805 ,21340 ,8879 ,17820 ,15104 ,7534 ,24323 ,21680 ,30302 ,18944 ,6536 ,23785 ,19221 ,2292 ,711 ,31344 ,13145 ,11972 ,18580 ,6289 ,22977 ,3580 ,15038 ,20710 ,12536 ,17728 ,12647 ,17284 ,12513 ,28917 ,14738 ,1992 ,10335 ,15231 ,14966 ,24930 ,30112 ,19584 ,25788 ,22556 ,3108 ,24218 ,15777 ,31112 ,20328 ,4164 ,22185 ,8973 ,1380 ,19516 ,25180 ,11797 ,3031 ,27548 ,23752 ,31439 ,23902 ,6256 ,15459 ,23935 ,22070 ,25709 ,17009 ,6722 ,8069 ,28745 ,14773 ,23685 ,31722 ,5645 ,5091 ,24747 ,26108 ,15849 ,27168 ,1092 ,9144 ,18070 ,
      1017 ,12438 ,26516 ,11299 ,3710 ,28778 ,3382 ,22856 ,14184 ,17872 ,5526 ,17519 ,24170 ,14329 ,21474 ,14028 ,27288 ,30638 ,18660 ,15978 ,12363 ,12936 ,8689 ,22338 ,7336 ,9674 ,19928 ,3758 ,12025 ,10046 ,177 ,6080 ,3466 ,3299 ,11015 ,19375 ,3259 ,5757 ,19593 ,24377 ,23279 ,14529 ,22687 ,1177 ,21288 ,8102 ,3750 ,17973 ,4309 ,23621 ,13011 ,29761 ,30147 ,31874 ,5145 ,22347 ,26662 ,9937 ,1648 ,4967 ,18827 ,20119 ,27963 ,10701 ,8006 ,20560 ,25076 ,27598 ,4269 ,25899 ,32383 ,7169 ,13726 ,15130 ,7232 ,18163 ,13661 ,31990 ,1969 ,883 ,4201 ,14564 ,23003 ,6410 ,22413 ,6755 ,8337 ,30138 ,3057 ,19877 ,9432 ,28536 ,14322 ,31748 ,19015 ,32225 ,26376 ,25365 ,25651 ,28826 ,10661 ,29670 ,9086 ,8764 ,25387 ,19257 ,17226 ,27651 ,19744 ,2822 ,15719 ,12854 ,26088 ,11423 ,2693 ,25500 ,3543 ,32467 ,30244 ,9843 ,2133 ,23543 ,1628 ,9412 ,1750 ,17042 ,31197 ,23443 ,9112 ,23870 ,30080 ,13113 ,18620 ,30270 ,32325 ,16238 ,11672 ,8579 ,32409 ,25220 ,25937 ,31755 ,10603 ,8363 ,28209 ,5171 ,15920 ,22904 ,19619 ,30380 ,26458 ,23612 ,16053 ,10752 ,23563 ,8715 ,6234 ,18443 ,3408 ,13273 ,18291 ,6327 ,20465 ,20596 ,10006 ,5678 ,14885 ,29138 ,619 ,29383 ,21118 ,18735 ,4760 ,6997 ,7328 ,30825 ,27931 ,22655 ,8657 ,26484 ,15687 ,1596 ,32351 ,22971 ,3376 ,32377 ,32319 ,20433 ,14911 ,4587 ,561 ,17611 ,21572 ,4443 ,32446 ,1575 ,24130 ,13075 ,20439 ,17799 ,29255 ,26716 ,28940 ,14249 ,10922 ,27363 ,14943 ,12781 ,9775 ,906 ,11152 ,6898 ,12804 ,16585 ,29112 ,13002 ,2187 ,31046 ,4619 ,28136 ,27493 ,14806 ,13494 ,20523 ,24016 ,21015 ,13413 ,21775 ,11259 ,6652 ,593 ,13830 ,22149 ,24518 ,1457 ,3430 ,7386 ,4034 ,7729 ,28334 ,2605 ,23314 ,17643 ,16856 ,24289 ,23718 ,6971 ,10523 ,2099 ,23245 ,2153 ,11638 ,31667 ,21176 ,30713 ,9554 ,
      3833 ,8248 ,12314 ,11210 ,8297 ,31578 ,14917 ,29294 ,11711 ,12225 ,29956 ,26564 ,9724 ,19022 ,16440 ,15283 ,5281 ,1212 ,29170 ,11505 ,6616 ,24780 ,14223 ,4958 ,30833 ,13765 ,17062 ,17981 ,30431 ,20802 ,26852 ,372 ,19452 ,4677 ,2940 ,6834 ,19837 ,27840 ,24104 ,9281 ,12672 ,2328 ,11750 ,22509 ,27006 ,15484 ,10038 ,20794 ,13552 ,5429 ,18358 ,20003 ,8482 ,4464 ,4417 ,12178 ,31701 ,25318 ,5710 ,9627 ,6950 ,5124 ,16538 ,24471 ,10185 ,19769 ,20628 ,15077 ,13686 ,15882 ,4593 ,32504 ,27801 ,32625 ,3942 ,21313 ,5873 ,8529 ,24195 ,28113 ,10947 ,24684 ,25566 ,6509 ,24621 ,7411 ,20497 ,26653 ,16730 ,11867 ,25962 ,21653 ,21467 ,10596 ,16433 ,4785 ,1493 ,2800 ,29890 ,27031 ,7129 ,28998 ,9749 ,8855 ,21210 ,5923 ,6359 ,13295 ,5898 ,26141 ,16929 ,7924 ,28060 ,4511 ,22262 ,11347 ,15001 ,27764 ,16559 ,16102 ,6180 ,28467 ,1770 ,26254 ,2658 ,11117 ,18323 ,21928 ,15577 ,5476 ,22789 ,12486 ,17186 ,28247 ,567 ,10801 ,8443 ,10251 ,27326 ,17701 ,22237 ,32232 ,4792 ,16635 ,31279 ,13903 ,21963 ,18553 ,5319 ,25812 ,21749 ,20110 ,30747 ,12100 ,7029 ,31317 ,22048 ,27201 ,7707 ,16907 ,8181 ,23162 ,21848 ,3081 ,29630 ,24816 ,7360 ,18920 ,19111 ,2211 ,10121 ,4137 ,16077 ,2458 ,169 ,26844 ,28662 ,22722 ,30857 ,14711 ,6001 ,1125 ,24492 ,16754 ,30771 ,21405 ,31217 ,24903 ,14122 ,13599 ,9050 ,24068 ,10446 ,4890 ,7847 ,3004 ,3503 ,18405 ,17617 ,762 ,9588 ,30942 ,29415 ,19489 ,6155 ,9177 ,20305 ,13471 ,30570 ,14630 ,4332 ,15432 ,24965 ,29825 ,10497 ,27954 ,13575 ,7474 ,23463 ,31412 ,1320 ,28685 ,651 ,1932 ,117 ,13968 ,18767 ,8042 ,9372 ,18103 ,2073 ,19197 ,26398 ,16178 ,15627 ,5618 ,11092 ,1515 ,2545 ,20955 ,16380 ,312 ,26946 ,5064 ,3882 ,21593 ,21150 ,28407 ,507 ,20050 ,29570 ,1065 ,7787 ,15372 ,57 ,252 ,
      237 ,7772 ,20035 ,29555 ,5049 ,16365 ,21578 ,21135 ,19182 ,9357 ,13953 ,18752 ,5603 ,26383 ,1500 ,2530 ,13456 ,6140 ,30927 ,29400 ,2989 ,10431 ,18390 ,17602 ,27939 ,24950 ,14615 ,4317 ,31397 ,13560 ,28670 ,636 ,16892 ,22033 ,12085 ,7014 ,18538 ,31264 ,25797 ,21734 ,10786 ,17171 ,5461 ,22774 ,17686 ,8428 ,32217 ,4777 ,26829 ,16062 ,2196 ,10106 ,3066 ,8166 ,24801 ,7345 ,16739 ,5986 ,22707 ,30842 ,24888 ,30756 ,13584 ,9035 ,24456 ,6935 ,25303 ,5695 ,19988 ,13537 ,4449 ,4402 ,9266 ,19822 ,4662 ,2925 ,22494 ,12657 ,15469 ,10023 ,15268 ,9709 ,12210 ,29941 ,11195 ,3818 ,31563 ,14902 ,4943 ,6601 ,1197 ,29155 ,17966 ,30818 ,20787 ,26837 ,4770 ,21452 ,11852 ,25947 ,6494 ,10932 ,7396 ,20482 ,32489 ,13671 ,19754 ,20613 ,21298 ,27786 ,8514 ,24180 ,7909 ,5883 ,5908 ,6344 ,27016 ,1478 ,28983 ,9734 ,16087 ,14986 ,4496 ,22247 ,26239 ,6165 ,11102 ,18308 ,23428 ,1735 ,23528 ,1613 ,25485 ,26073 ,32452 ,30229 ,8749 ,10646 ,25350 ,25636 ,27636 ,25372 ,2807 ,15704 ,868 ,13646 ,15115 ,7217 ,27583 ,7991 ,25884 ,32368 ,30123 ,22398 ,14549 ,22988 ,28521 ,3042 ,31733 ,19000 ,6065 ,12010 ,9659 ,19913 ,15963 ,27273 ,12921 ,8674 ,22841 ,3695 ,12423 ,26501 ,17504 ,14169 ,14314 ,21459 ,17958 ,21273 ,14514 ,22672 ,19360 ,3451 ,5742 ,19578 ,22332 ,30132 ,23606 ,12996 ,4952 ,26647 ,20104 ,27948 ,17596 ,14896 ,32362 ,32304 ,26469 ,27916 ,1581 ,32336 ,29123 ,9991 ,6312 ,20450 ,18720 ,604 ,6982 ,7313 ,8348 ,25922 ,8564 ,32394 ,13098 ,9097 ,30255 ,32310 ,23597 ,19604 ,5156 ,15905 ,8700 ,16038 ,18428 ,3393 ,20508 ,27478 ,31031 ,4604 ,6883 ,9760 ,16570 ,29097 ,17784 ,24115 ,4428 ,32431 ,14234 ,29240 ,27348 ,14928 ,28319 ,7371 ,24503 ,1442 ,21760 ,24001 ,6637 ,578 ,10508 ,24274 ,23299 ,17628 ,11623 ,2084 ,21161 ,30698 ,
      11058 ,14088 ,5839 ,30397 ,4726 ,31633 ,24136 ,14288 ,25259 ,16801 ,12613 ,25124 ,17922 ,25658 ,29897 ,19636 ,21534 ,3793 ,9313 ,23073 ,27895 ,16344 ,17558 ,26475 ,22663 ,18202 ,8122 ,23629 ,18494 ,5437 ,22730 ,32136 ,2763 ,8936 ,1691 ,14389 ,824 ,21352 ,18956 ,15937 ,14470 ,13358 ,26603 ,22921 ,17460 ,28006 ,19869 ,11859 ,6593 ,15243 ,24230 ,5188 ,17740 ,24539 ,29053 ,11984 ,6268 ,10355 ,27872 ,19528 ,13054 ,28757 ,15861 ,28226 ,11606 ,28302 ,6866 ,17767 ,18703 ,17579 ,13081 ,23580 ,28504 ,851 ,25468 ,8732 ,17487 ,6048 ,19343 ,22315 ,24871 ,26812 ,18521 ,10769 ,5586 ,220 ,2972 ,27922 ,17949 ,15251 ,19971 ,9249 ,21281 ,4753 ,26999 ,16070 ,17679 ,17497 ,17453 ,18460 ,17470 ,11589 ,5569 ,17932 ,18477 ,21517 ,4709 ,25242 ,17443 ,2746 ,17723 ,6251 ,17514 ,1172 ,18158 ,27646 ,25215 ,18730 ,14244 ,3425 ,26559 ,22504 ,21308 ,13290 ,17696 ,4132 ,19484 ,5613 ,18747 ,22769 ,2920 ,20608 ,25631 ,26496 ,20445 ,32426 ,25119 ,22916 ,8727 ,25237 ,25232 ,28833 ,27038 ,13125 ,12743 ,6910 ,28148 ,8596 ,14261 ,31136 ,7275 ,1587 ,3442 ,2012 ,15516 ,21787 ,5812 ,16868 ,11650 ,11689 ,32057 ,6422 ,28548 ,31772 ,18175 ,19058 ,10070 ,27610 ,27663 ,14830 ,9475 ,28838 ,18467 ,25512 ,9424 ,25954 ,1189 ,19963 ,20826 ,19387 ,23046 ,29773 ,4979 ,10620 ,27225 ,15990 ,3770 ,8380 ,17531 ,28709 ,29725 ,11311 ,2277 ,6521 ,21665 ,30287 ,21325 ,30904 ,17805 ,15089 ,13307 ,30325 ,2360 ,27043 ,2736 ,11359 ,26266 ,18637 ,22521 ,2900 ,1671 ,6846 ,11832 ,20015 ,9639 ,32342 ,5733 ,11517 ,17993 ,16255 ,26576 ,31240 ,12704 ,11222 ,4149 ,15762 ,22541 ,3093 ,15216 ,14723 ,24915 ,30097 ,3565 ,18565 ,31329 ,13130 ,17713 ,15023 ,17269 ,12498 ,25694 ,15444 ,31424 ,23887 ,19501 ,22170 ,11782 ,3016 ,5630 ,14758 ,6707 ,8054 ,15834 ,5076 ,1077 ,9129 ,
      28374 ,1899 ,18887 ,16602 ,26620 ,21895 ,29261 ,20761 ,22938 ,13240 ,13797 ,12748 ,22305 ,10668 ,7136 ,12821 ,13375 ,8403 ,1813 ,20179 ,19551 ,18037 ,30993 ,29129 ,8665 ,26204 ,5777 ,13019 ,14487 ,18366 ,30865 ,31501 ,28023 ,16972 ,18013 ,28572 ,3668 ,1879 ,22565 ,11169 ,27458 ,1715 ,22013 ,6915 ,17477 ,14068 ,6402 ,6501 ,29933 ,10761 ,31055 ,923 ,19886 ,4055 ,17094 ,9683 ,11876 ,3128 ,12590 ,13774 ,12894 ,12109 ,7483 ,9792 ,21369 ,23209 ,16275 ,15178 ,7964 ,9334 ,26722 ,4636 ,20671 ,32570 ,7563 ,28153 ,841 ,10838 ,30463 ,17849 ,29477 ,21709 ,32660 ,31063 ,18973 ,15323 ,3985 ,9997 ,15954 ,24238 ,20834 ,23814 ,14522 ,29376 ,2321 ,2204 ,17164 ,3688 ,13351 ,14823 ,1708 ,16476 ,26884 ,24430 ,14406 ,16675 ,26005 ,8601 ,25458 ,2404 ,10273 ,27510 ,8953 ,12060 ,404 ,26310 ,25609 ,5027 ,29191 ,13511 ,20995 ,23850 ,3279 ,20540 ,2780 ,8228 ,23142 ,4870 ,24556 ,30010 ,11537 ,17313 ,29213 ,23094 ,28946 ,28957 ,25749 ,20739 ,30207 ,14266 ,17757 ,29677 ,29005 ,19295 ,3996 ,5961 ,3609 ,26733 ,29070 ,26895 ,29202 ,6318 ,12001 ,22576 ,17105 ,31934 ,31004 ,31373 ,16216 ,29272 ,23350 ,22585 ,31477 ,27380 ,24247 ,20252 ,29999 ,26213 ,5205 ,16483 ,1244 ,31141 ,11596 ,7653 ,4193 ,10939 ,15260 ,24863 ,29469 ,18211 ,1415 ,2021 ,11526 ,14960 ,12357 ,22407 ,19613 ,12798 ,6610 ,24615 ,5313 ,24959 ,2983 ,11189 ,27577 ,13092 ,27889 ,5580 ,14255 ,11826 ,19545 ,18967 ,29064 ,7280 ,17569 ,9002 ,4369 ,24147 ,10372 ,10081 ,4990 ,23964 ,7286 ,457 ,25738 ,20456 ,9650 ,31468 ,24397 ,17816 ,6285 ,24926 ,11793 ,23681 ,28774 ,12932 ,5753 ,31870 ,25895 ,6751 ,29666 ,32463 ,30266 ,30376 ,5674 ,1592 ,13071 ,16581 ,6648 ,23714 ,31574 ,24776 ,27836 ,4460 ,15878 ,7407 ,28994 ,27760 ,28243 ,25808 ,24812 ,1121 ,18401 ,29821 ,18099 ,21589 ,
      16361 ,10427 ,31260 ,8162 ,13533 ,3814 ,10928 ,1474 ,26069 ,7987 ,27269 ,3447 ,27912 ,9093 ,9756 ,23997 ,31629 ,16340 ,21348 ,24535 ,17575 ,216 ,11585 ,18726 ,26492 ,31132 ,19054 ,29769 ,30900 ,20011 ,14719 ,22166 ,21891 ,18033 ,1875 ,4051 ,9330 ,15319 ,16472 ,5023 ,23090 ,26891 ,20248 ,2017 ,5576 ,453 ,6747 ,7403 ,3810 ,212 ,15315 ,32738 ,29528 ,32742 ,1233 ,7746 ,690 ,20870 ,11035 ,28351 ,21551 ,996 ,10164 ,15556 ,20367 ,28592 ,11448 ,6669 ,8139 ,29532 ,27369 ,14589 ,23646 ,4835 ,12257 ,15521 ,26802 ,30663 ,32101 ,11276 ,18219 ,2505 ,5372 ,931 ,9008 ,32746 ,23339 ,610 ,22832 ,5196 ,19395 ,13847 ,22680 ,21111 ,11743 ,10114 ,5454 ,12416 ,26596 ,9468 ,22006 ,1237 ,20241 ,13430 ,9865 ,30515 ,4536 ,21792 ,18511 ,16124 ,17361 ,24709 ,19672 ,13928 ,27707 ,21032 ,22747 ,7750 ,29988 ,10405 ,32153 ,15797 ,7072 ,14655 ,32190 ,9519 ,337 ,24033 ,27151 ,16992 ,25163 ,23735 ,12630 ,694 ,14949 ,25771 ,25141 ,18865 ,23506 ,5817 ,9239 ,8771 ,8862 ,24306 ,16818 ,6115 ,29326 ,27082 ,4375 ,20874 ,1404 ,6988 ,14160 ,7644 ,3319 ,10540 ,25276 ,19158 ,30058 ,12292 ,25675 ,2258 ,12724 ,32038 ,6574 ,11039 ,24852 ,17660 ,7890 ,24437 ,13437 ,16873 ,17939 ,23409 ,8329 ,20489 ,31555 ,2964 ,3977 ,23331 ,29914 ,28355 ,29458 ,17145 ,19653 ,20348 ,31610 ,21872 ,31536 ,27132 ,18791 ,2622 ,31650 ,2588 ,11242 ,22132 ,10905 ,21555 ,12787 ,2170 ,6217 ,28192 ,18603 ,11655 ,4743 ,18274 ,15670 ,3359 ,18810 ,4292 ,3242 ,23262 ,24153 ,1000 ,12346 ,7319 ,14305 ,4184 ,4252 ,13709 ,19727 ,26359 ,3526 ,2116 ,2641 ,28043 ,7112 ,21193 ,5856 ,10168 ,24604 ,16713 ,30414 ,5264 ,8280 ,11694 ,26989 ,19435 ,8465 ,31684 ,14105 ,28645 ,29613 ,19094 ,22220 ,15560 ,5302 ,30730 ,1303 ,30553 ,3486 ,9571 ,11075 ,100 ,3865 ,490 ,
      20893 ,4075 ,8793 ,6772 ,9492 ,20371 ,9781 ,29699 ,28855 ,17386 ,3151 ,32062 ,32126 ,25394 ,21217 ,22430 ,14847 ,16013 ,8887 ,2851 ,10378 ,28596 ,12883 ,8354 ,15695 ,19286 ,31894 ,30155 ,27680 ,8490 ,6009 ,27404 ,25529 ,10298 ,2380 ,31796 ,30488 ,11452 ,3117 ,23020 ,13188 ,14413 ,9872 ,6427 ,18484 ,3205 ,7161 ,32496 ,4394 ,23572 ,4628 ,14581 ,9441 ,6673 ,12579 ,19937 ,25971 ,12556 ,29030 ,17071 ,20214 ,7038 ,23472 ,4218 ,19075 ,22113 ,27063 ,32019 ,32719 ,8143 ,912 ,9449 ,26291 ,15159 ,20160 ,28553 ,18192 ,17294 ,23945 ,31851 ,1423 ,32285 ,7198 ,19894 ,10087 ,29536 ,29922 ,25928 ,27627 ,17748 ,23054 ,14370 ,19368 ,20589 ,6827 ,3074 ,7007 ,19906 ,14382 ,31765 ,28565 ,27373 ,4044 ,32031 ,31789 ,32000 ,2832 ,31777 ,8112 ,31820 ,32254 ,14339 ,6439 ,8539 ,26151 ,31808 ,15494 ,14593 ,17083 ,19032 ,2468 ,2863 ,30167 ,32242 ,32074 ,9187 ,1525 ,6784 ,29790 ,27729 ,30345 ,31839 ,426 ,23650 ,11158 ,7249 ,7622 ,26182 ,22376 ,18180 ,23063 ,19264 ,5930 ,31903 ,29345 ,9966 ,32539 ,15147 ,4996 ,4839 ,3657 ,8570 ,10637 ,20730 ,26173 ,20148 ,1848 ,6470 ,10730 ,13743 ,27101 ,17114 ,24406 ,32007 ,20843 ,12261 ,16961 ,5786 ,19404 ,16682 ,30522 ,19063 ,21524 ,3328 ,4261 ,13678 ,19980 ,18695 ,7956 ,8131 ,32711 ,15525 ,18002 ,1986 ,30632 ,14558 ,5165 ,900 ,1206 ,24678 ,13897 ,14624 ,6134 ,9703 ,13640 ,25916 ,3787 ,26806 ,6904 ,2894 ,8397 ,21703 ,5955 ,10075 ,16334 ,2499 ,6109 ,4286 ,16007 ,32279 ,9960 ,32273 ,23970 ,30667 ,27447 ,32400 ,25341 ,30198 ,22367 ,7186 ,27242 ,21428 ,21242 ,12965 ,28726 ,11953 ,13327 ,14358 ,16313 ,32105 ,14057 ,25093 ,2715 ,17901 ,22473 ,27615 ,17548 ,22284 ,26781 ,9218 ,16837 ,1556 ,22885 ,20577 ,29742 ,11280 ,6391 ,28807 ,11328 ,15058 ,11486 ,6815 ,14692 ,12467 ,15413 ,8023 ,
      31153 ,21054 ,11379 ,27392 ,26332 ,18223 ,12810 ,17243 ,25032 ,26745 ,31946 ,27668 ,14278 ,17233 ,6366 ,17325 ,3338 ,23976 ,17828 ,19274 ,7292 ,2509 ,22294 ,13104 ,1604 ,17304 ,31830 ,31882 ,3215 ,4472 ,1133 ,25404 ,10559 ,31075 ,23826 ,2839 ,28165 ,5376 ,13229 ,15190 ,8613 ,26012 ,4543 ,14835 ,4716 ,26322 ,20552 ,19761 ,6927 ,28294 ,23201 ,28584 ,22105 ,935 ,13786 ,15736 ,28896 ,20191 ,13031 ,12871 ,12760 ,14007 ,28092 ,16614 ,7663 ,943 ,13859 ,29687 ,15533 ,9012 ,16591 ,6681 ,21804 ,10848 ,2414 ,9480 ,14078 ,21044 ,14667 ,10678 ,2029 ,30673 ,16134 ,4063 ,463 ,32750 ,28363 ,9103 ,23419 ,24547 ,29781 ,8781 ,3459 ,18284 ,19445 ,8174 ,16885 ,6058 ,2756 ,32050 ,28016 ,23343 ,21884 ,25668 ,25522 ,27094 ,10552 ,28843 ,5829 ,11369 ,15033 ,23747 ,14179 ,23274 ,13721 ,25382 ,11667 ,614 ,29250 ,22144 ,11706 ,12667 ,27796 ,21205 ,8438 ,19106 ,9583 ,26393 ,19177 ,10781 ,9261 ,32484 ,8744 ,22836 ,29118 ,17779 ,25254 ,14465 ,28499 ,18472 ,25114 ,27658 ,13302 ,3560 ,22933 ,27453 ,20666 ,14401 ,25744 ,5200 ,19540 ,30261 ,26064 ,23085 ,23641 ,9860 ,25136 ,7885 ,6212 ,30409 ,28850 ,13183 ,26286 ,31784 ,7617 ,19399 ,8392 ,2710 ,25027 ,8608 ,21799 ,25517 ,25249 ,25022 ,25068 ,20620 ,25295 ,6858 ,16267 ,11440 ,27055 ,13851 ,1802 ,30299 ,13142 ,12533 ,10332 ,3105 ,1377 ,23899 ,8066 ,26105 ,26513 ,5523 ,18657 ,19925 ,11012 ,22684 ,13008 ,1645 ,25073 ,7229 ,23000 ,9429 ,25648 ,17223 ,2690 ,1625 ,30077 ,32406 ,15917 ,23560 ,20462 ,21115 ,8654 ,32316 ,32443 ,28937 ,11149 ,4616 ,13410 ,1454 ,17640 ,2150 ,12311 ,29953 ,29167 ,17059 ,2937 ,11747 ,18355 ,5707 ,20625 ,3939 ,25563 ,25959 ,29887 ,6356 ,22259 ,1767 ,22786 ,27323 ,21960 ,7026 ,21845 ,10118 ,30854 ,31214 ,7844 ,29412 ,4329 ,23460 ,18764 ,15624 ,26943 ,29567 ,
      20032 ,13950 ,30924 ,14612 ,12082 ,5458 ,2193 ,22704 ,25300 ,4659 ,12207 ,1194 ,11849 ,19751 ,5905 ,4493 ,23525 ,25347 ,15112 ,14546 ,9656 ,12420 ,14511 ,23603 ,32359 ,6309 ,8561 ,5153 ,31028 ,4425 ,24500 ,23296 ,5836 ,12610 ,9310 ,8119 ,1688 ,26600 ,24227 ,27869 ,6863 ,25465 ,18518 ,19968 ,17450 ,4706 ,18155 ,21305 ,2917 ,8724 ,28145 ,15513 ,28545 ,9472 ,20823 ,3767 ,21662 ,2357 ,1668 ,17990 ,22538 ,31326 ,31421 ,6704 ,18884 ,13794 ,1810 ,5774 ,18010 ,22010 ,31052 ,12587 ,16272 ,7560 ,32657 ,20831 ,13348 ,26002 ,401 ,3276 ,11534 ,30204 ,3606 ,17102 ,31474 ,1241 ,29466 ,19610 ,27574 ,29061 ,4987 ,24394 ,5750 ,5671 ,27833 ,24809 ,31257 ,27266 ,21345 ,19051 ,1872 ,20245 ,15312 ,11032 ,11445 ,12254 ,5369 ,19392 ,26593 ,4533 ,27704 ,7069 ,25160 ,23503 ,29323 ,3316 ,12721 ,13434 ,3974 ,31607 ,11239 ,18600 ,3239 ,4249 ,7109 ,8277 ,29610 ,3483 ,8790 ,3148 ,8884 ,31891 ,2377 ,9869 ,4625 ,29027 ,27060 ,20157 ,7195 ,23051 ,14379 ,2829 ,26148 ,30164 ,30342 ,22373 ,32536 ,26170 ,24403 ,30519 ,7953 ,5162 ,13637 ,5952 ,9957 ,22364 ,13324 ,22470 ,22882 ,11483 ,11376 ,31943 ,17825 ,31827 ,23823 ,4540 ,23198 ,13028 ,13856 ,2411 ,16131 ,29778 ,2753 ,10549 ,13718 ,27793 ,9258 ,28496 ,20663 ,23638 ,26283 ,21796 ,16264 ,10329 ,18654 ,22997 ,15914 ,11146 ,29164 ,25560 ,21957 ,4326 ,30921 ,12204 ,15109 ,8558 ,9307 ,18515 ,28142 ,1665 ,1807 ,32654 ,3603 ,4984 ,21342 ,5366 ,29320 ,3236 ,8881 ,7192 ,32533 ,9954 ,17822 ,16128 ,20660 ,15911 ,15106 ,3600 ,32530 ,32527 ,7536 ,19798 ,785 ,26679 ,24325 ,11896 ,7539 ,20136 ,21682 ,17365 ,10827 ,14444 ,30304 ,16780 ,19801 ,10625 ,18946 ,13219 ,4814 ,18844 ,6538 ,25859 ,788 ,6458 ,23787 ,24713 ,30452 ,27980 ,19223 ,9903 ,26682 ,10718 ,2294 ,28433 ,10217 ,7440 ,
      713 ,12129 ,24328 ,12953 ,31346 ,19676 ,27499 ,19317 ,13147 ,11917 ,11899 ,27230 ,11974 ,15726 ,16936 ,12380 ,18582 ,27248 ,7542 ,30186 ,6291 ,13932 ,25447 ,8706 ,22979 ,31925 ,20139 ,22355 ,3582 ,12186 ,16762 ,25841 ,15040 ,11935 ,21685 ,32261 ,20712 ,27711 ,16664 ,18677 ,12538 ,10280 ,17368 ,15995 ,17730 ,22095 ,31982 ,8521 ,12649 ,6040 ,10830 ,30655 ,17286 ,21036 ,25994 ,28276 ,12515 ,13165 ,14447 ,27435 ,28919 ,5505 ,3921 ,27305 ,14740 ,15744 ,30307 ,2882 ,1994 ,22751 ,14812 ,19945 ,10337 ,8918 ,16783 ,3775 ,15233 ,28284 ,21499 ,1154 ,14968 ,21434 ,19804 ,9691 ,24932 ,7754 ,17153 ,16044 ,30114 ,11992 ,10628 ,13628 ,19586 ,14878 ,24097 ,7353 ,25790 ,12914 ,18949 ,10063 ,22558 ,29992 ,16465 ,24845 ,3110 ,16954 ,13222 ,8385 ,24220 ,23191 ,16657 ,12042 ,15779 ,12398 ,4817 ,2487 ,31114 ,10409 ,26873 ,194 ,20330 ,2240 ,18847 ,6097 ,4166 ,2570 ,5246 ,28627 ,22187 ,19694 ,6541 ,9206 ,8975 ,32157 ,13500 ,5543 ,1382 ,30971 ,25862 ,17536 ,19518 ,12861 ,7931 ,25425 ,25182 ,21248 ,791 ,17889 ,11799 ,15801 ,25598 ,18434 ,3033 ,31364 ,6461 ,22461 ,27550 ,4919 ,26436 ,14201 ,23754 ,7503 ,23790 ,14346 ,31441 ,7076 ,12049 ,17417 ,23904 ,27517 ,24716 ,28714 ,6258 ,28886 ,1961 ,24187 ,15461 ,19335 ,30455 ,32093 ,23937 ,14659 ,393 ,21491 ,22072 ,3182 ,27983 ,14045 ,25711 ,1344 ,10979 ,29854 ,17011 ,9812 ,19226 ,28795 ,6724 ,32194 ,20529 ,18132 ,8071 ,24346 ,9906 ,29730 ,28747 ,13997 ,30607 ,3727 ,14775 ,12971 ,26685 ,1544 ,23687 ,9523 ,20984 ,3399 ,31724 ,16207 ,10721 ,22873 ,5647 ,30794 ,22624 ,20402 ,5093 ,12147 ,2297 ,6803 ,24749 ,341 ,8217 ,26533 ,26110 ,8824 ,28436 ,11316 ,15851 ,28082 ,24653 ,21622 ,27170 ,20079 ,10220 ,12455 ,1094 ,24037 ,23131 ,4106 ,9146 ,731 ,7443 ,15401 ,18072 ,20924 ,281 ,1034 ,
      1019 ,18057 ,716 ,7428 ,12440 ,27155 ,24022 ,23116 ,26518 ,24734 ,12132 ,2282 ,11301 ,26095 ,28067 ,24638 ,3712 ,28732 ,24331 ,9891 ,28780 ,16996 ,32179 ,20514 ,3384 ,23672 ,12956 ,26670 ,22858 ,31709 ,30779 ,22609 ,14186 ,27535 ,31349 ,6446 ,17874 ,25167 ,15786 ,25583 ,5528 ,8960 ,19679 ,6526 ,17521 ,1367 ,12846 ,7916 ,24172 ,6243 ,27502 ,24701 ,14331 ,23739 ,7061 ,12034 ,21476 ,23922 ,19320 ,30440 ,14030 ,22057 ,1329 ,10964 ,27290 ,28904 ,13150 ,14432 ,30640 ,12634 ,21021 ,25979 ,18662 ,20697 ,11920 ,21670 ,15980 ,12523 ,22080 ,31967 ,12365 ,11959 ,11902 ,11884 ,12938 ,698 ,19661 ,27484 ,8691 ,6276 ,27233 ,7527 ,22340 ,22964 ,12171 ,16747 ,7338 ,19571 ,11977 ,10613 ,9676 ,14953 ,7739 ,17138 ,19930 ,1979 ,15729 ,30292 ,3760 ,10322 ,28269 ,21484 ,12027 ,24205 ,16939 ,13207 ,10048 ,25775 ,29977 ,16450 ,179 ,31099 ,12383 ,4802 ,6082 ,20315 ,2555 ,5231 ,3468 ,7094 ,18585 ,3224 ,3301 ,25145 ,13419 ,3959 ,11017 ,1857 ,27251 ,21330 ,19377 ,11430 ,4518 ,27689 ,3261 ,13333 ,7545 ,32642 ,5759 ,18869 ,21995 ,31037 ,19595 ,31459 ,30189 ,3591 ,24379 ,27559 ,5656 ,27818 ,23281 ,31013 ,6294 ,8546 ,14531 ,23510 ,12405 ,14496 ,22689 ,12067 ,13935 ,30909 ,1179 ,25285 ,19736 ,5890 ,21290 ,17435 ,25450 ,18503 ,8104 ,5821 ,26585 ,24212 ,3752 ,28530 ,8709 ,28130 ,17975 ,21647 ,31311 ,31406 ,4311 ,29149 ,22982 ,15899 ,23623 ,9243 ,21781 ,16249 ,13013 ,23808 ,31928 ,17810 ,29763 ,13841 ,10534 ,13703 ,30149 ,14364 ,20142 ,7180 ,31876 ,8775 ,9854 ,4610 ,5147 ,24388 ,22358 ,32521 ,22349 ,13622 ,22455 ,22867 ,26664 ,7521 ,3585 ,32515 ,9939 ,8866 ,16113 ,20645 ,1650 ,9292 ,12189 ,15094 ,4969 ,1792 ,5351 ,29305 ,18829 ,18931 ,16765 ,19786 ,20121 ,24310 ,17350 ,10812 ,27965 ,23772 ,25844 ,773 ,10703 ,19208 ,28418 ,10202 ,
      8008 ,14677 ,15043 ,11471 ,20562 ,16822 ,11265 ,6376 ,25078 ,16298 ,11938 ,13312 ,27600 ,2700 ,22269 ,26766 ,4271 ,16319 ,21688 ,5940 ,25901 ,6119 ,26791 ,6889 ,32385 ,23955 ,32264 ,9945 ,7171 ,25326 ,21413 ,21227 ,13728 ,1833 ,20715 ,26158 ,15132 ,29330 ,4824 ,3642 ,7234 ,411 ,27714 ,30330 ,18165 ,7607 ,19249 ,5915 ,13663 ,21509 ,16667 ,30507 ,31992 ,27086 ,12246 ,16946 ,1971 ,32696 ,18680 ,7941 ,885 ,30617 ,24663 ,13882 ,4203 ,20199 ,12541 ,29015 ,14566 ,4379 ,6658 ,12564 ,23005 ,30473 ,10283 ,2365 ,6412 ,13173 ,3190 ,7146 ,22415 ,32111 ,17371 ,3136 ,6757 ,20878 ,20356 ,9766 ,8339 ,10363 ,15998 ,8872 ,30140 ,15680 ,8475 ,5994 ,3059 ,19353 ,17733 ,23039 ,19879 ,1408 ,29521 ,29907 ,9434 ,32704 ,22098 ,27048 ,28538 ,26276 ,17279 ,23930 ,14324 ,8097 ,31985 ,2817 ,31750 ,6992 ,27358 ,4029 ,19017 ,15479 ,8524 ,26136 ,32227 ,2453 ,9172 ,1510 ,26378 ,8423 ,12652 ,27781 ,25367 ,14164 ,599 ,29235 ,25653 ,28001 ,6043 ,2741 ,28828 ,25507 ,11354 ,15018 ,10663 ,14063 ,10833 ,2399 ,29672 ,7648 ,8997 ,16576 ,9088 ,448 ,30658 ,16119 ,8766 ,23404 ,18269 ,19430 ,25389 ,3200 ,17289 ,31815 ,19259 ,3323 ,2494 ,22279 ,17228 ,26317 ,21039 ,11364 ,27653 ,25017 ,17218 ,6351 ,19746 ,4701 ,25997 ,4528 ,2824 ,10544 ,5361 ,13214 ,15721 ,22090 ,28279 ,23186 ,12856 ,28881 ,13992 ,28077 ,26090 ,1362 ,12518 ,10317 ,11425 ,25280 ,13836 ,1787 ,2695 ,7602 ,13168 ,26271 ,25502 ,25012 ,25007 ,25053 ,3545 ,25099 ,14450 ,28484 ,32469 ,19162 ,22821 ,29103 ,30246 ,25729 ,27438 ,20651 ,9845 ,26049 ,7870 ,6197 ,2135 ,13395 ,28922 ,11134 ,23545 ,30062 ,21100 ,8639 ,1630 ,10997 ,5508 ,18642 ,9414 ,25058 ,17208 ,2675 ,1752 ,29872 ,3924 ,25548 ,17044 ,12296 ,11732 ,18340 ,31199 ,21830 ,27308 ,21945 ,23445 ,7829 ,15609 ,26928 ,
      9114 ,15819 ,14743 ,6692 ,23872 ,25679 ,22155 ,11767 ,30082 ,15201 ,15747 ,22526 ,13115 ,3550 ,15008 ,17254 ,18622 ,2721 ,30310 ,2345 ,30272 ,2262 ,30889 ,17790 ,32327 ,11817 ,2885 ,1656 ,16240 ,5718 ,31225 ,12689 ,11674 ,5797 ,1997 ,15501 ,8581 ,12728 ,31121 ,7260 ,32411 ,25616 ,22754 ,2905 ,25222 ,25104 ,28818 ,27023 ,25939 ,18452 ,14815 ,9460 ,31757 ,32042 ,19043 ,10055 ,10605 ,23031 ,19948 ,20811 ,8365 ,27210 ,28694 ,29710 ,28211 ,13039 ,10340 ,27857 ,5173 ,6578 ,24524 ,29038 ,15922 ,809 ,8921 ,1676 ,22906 ,14455 ,27991 ,19854 ,19621 ,17907 ,16786 ,12598 ,30382 ,11043 ,31618 ,24121 ,26460 ,27880 ,3778 ,9298 ,23614 ,22648 ,5422 ,22715 ,16055 ,21266 ,15236 ,19956 ,10754 ,24856 ,205 ,2957 ,23565 ,18688 ,28287 ,6851 ,8717 ,28489 ,6033 ,19328 ,6236 ,17428 ,21502 ,4694 ,18445 ,17664 ,11574 ,5554 ,3410 ,25200 ,1157 ,18143 ,13275 ,26544 ,4117 ,19469 ,18293 ,26224 ,14971 ,4481 ,6329 ,7894 ,1463 ,28968 ,20467 ,6479 ,21437 ,11837 ,20598 ,32474 ,27771 ,8499 ,10008 ,22479 ,19807 ,4647 ,5680 ,24441 ,13522 ,4434 ,14887 ,11180 ,9694 ,12195 ,29140 ,4928 ,30803 ,20772 ,621 ,31382 ,24935 ,14600 ,29385 ,13441 ,10416 ,18375 ,21120 ,5034 ,7757 ,20020 ,18737 ,19167 ,26368 ,1485 ,4762 ,17671 ,17156 ,5446 ,6999 ,16877 ,31249 ,25782 ,7330 ,3051 ,16047 ,2181 ,30827 ,16724 ,30741 ,13569 ,27933 ,4937 ,30117 ,23591 ,22657 ,17943 ,3436 ,5727 ,8659 ,15948 ,11995 ,9644 ,26486 ,22826 ,14154 ,14299 ,15689 ,27621 ,10631 ,25335 ,1598 ,23413 ,26058 ,32437 ,32353 ,27568 ,13631 ,15100 ,22973 ,30108 ,3027 ,31718 ,3378 ,8685 ,19589 ,5141 ,32379 ,8333 ,9082 ,30240 ,32321 ,26454 ,14881 ,32347 ,20435 ,29108 ,589 ,6967 ,14913 ,14219 ,24100 ,4413 ,4589 ,20493 ,9745 ,16555 ,563 ,21745 ,7356 ,24488 ,17613 ,10493 ,2069 ,21146 ,
      21574 ,18386 ,25793 ,24797 ,4445 ,31559 ,7392 ,28979 ,32448 ,25880 ,12917 ,5738 ,1577 ,30251 ,16566 ,6633 ,24132 ,17554 ,18952 ,29049 ,13077 ,2968 ,5565 ,14240 ,20441 ,7271 ,10066 ,4975 ,17801 ,9635 ,24911 ,11778 ,29257 ,30989 ,22561 ,17090 ,26718 ,3981 ,26880 ,29187 ,28942 ,29198 ,29995 ,11522 ,14251 ,25734 ,29662 ,28990 ,10924 ,11581 ,16468 ,1229 ,27365 ,23335 ,20237 ,29984 ,14945 ,1400 ,24848 ,29454 ,12783 ,12342 ,24600 ,5298 ,9777 ,12879 ,3113 ,12575 ,908 ,29918 ,4040 ,17079 ,11154 ,3653 ,16957 ,17998 ,6900 ,27443 ,14053 ,6387 ,12806 ,22290 ,13225 ,13782 ,16587 ,28359 ,21880 ,29246 ,29114 ,19536 ,8388 ,1798 ,13004 ,8650 ,18351 ,30850 ,2189 ,14507 ,24223 ,20819 ,31048 ,29462 ,15308 ,3970 ,4621 ,7949 ,23194 ,16260 ,28138 ,20656 ,10823 ,30448 ,27495 ,25443 ,16660 ,25990 ,14808 ,17149 ,16461 ,26869 ,13496 ,25594 ,12045 ,389 ,20525 ,20980 ,8213 ,23127 ,24018 ,32175 ,15782 ,7057 ,21017 ,19657 ,7735 ,29973 ,13415 ,21991 ,12401 ,26581 ,21777 ,9850 ,16109 ,17346 ,11261 ,26787 ,4820 ,12242 ,6654 ,20352 ,29517 ,27354 ,595 ,8993 ,2490 ,5357 ,13832 ,22817 ,21096 ,11728 ,22151 ,30885 ,31117 ,19039 ,24520 ,31614 ,201 ,11570 ,1459 ,13518 ,10412 ,31245 ,3432 ,26054 ,9078 ,9741 ,7388 ,5561 ,26876 ,20233 ,4036 ,21876 ,15304 ,16457 ,7731 ,29513 ,197 ,15300 ,28336 ,675 ,981 ,10149 ,2607 ,31521 ,20333 ,31595 ,23316 ,31540 ,28340 ,29443 ,17645 ,6559 ,2243 ,12709 ,16858 ,7875 ,23394 ,8314 ,24291 ,9224 ,18850 ,23491 ,23720 ,27136 ,679 ,14934 ,6973 ,4360 ,6100 ,29311 ,10525 ,14145 ,19143 ,30043 ,2101 ,19712 ,4169 ,4237 ,23247 ,18795 ,985 ,12331 ,2155 ,10890 ,2573 ,11227 ,11640 ,6202 ,18259 ,15655 ,31669 ,26974 ,5249 ,8265 ,21178 ,2626 ,10153 ,24589 ,30715 ,22205 ,28630 ,29598 ,9556 ,1288 ,85 ,3850 ,
      3835 ,9541 ,22190 ,28615 ,8250 ,31654 ,2611 ,10138 ,12316 ,23232 ,19697 ,4154 ,11212 ,2140 ,6187 ,18244 ,8299 ,16843 ,6544 ,2228 ,31580 ,2592 ,31525 ,28325 ,14919 ,23705 ,9209 ,18835 ,29296 ,6958 ,14130 ,19128 ,11713 ,13817 ,8978 ,2475 ,12227 ,11246 ,20337 ,29502 ,29958 ,21002 ,32160 ,15767 ,26566 ,13400 ,9835 ,16094 ,9726 ,3417 ,13503 ,10397 ,19024 ,22136 ,31599 ,186 ,16442 ,4021 ,5546 ,26861 ,15285 ,7716 ,660 ,966 ,5283 ,12768 ,1385 ,24833 ,1214 ,10909 ,23320 ,20222 ,29172 ,26703 ,30974 ,22546 ,11507 ,28927 ,25719 ,29647 ,6618 ,1562 ,25865 ,12902 ,24782 ,21559 ,31544 ,7377 ,14225 ,13062 ,17539 ,18937 ,4960 ,20426 ,9620 ,24896 ,30835 ,12989 ,19521 ,8373 ,13767 ,12791 ,28344 ,21865 ,17064 ,893 ,12864 ,3098 ,17983 ,11139 ,27428 ,14038 ,30433 ,28123 ,7934 ,23179 ,20804 ,2174 ,29447 ,15293 ,26854 ,14793 ,25428 ,16645 ,374 ,13481 ,20965 ,8198 ,19454 ,13260 ,25185 ,1142 ,4679 ,6221 ,17649 ,11559 ,2942 ,10739 ,21251 ,15221 ,6836 ,23550 ,28474 ,6018 ,19839 ,22891 ,794 ,8906 ,27842 ,28196 ,6563 ,24509 ,24106 ,30367 ,17892 ,16771 ,9283 ,26445 ,22633 ,5407 ,12674 ,16225 ,11802 ,2870 ,2330 ,18607 ,2247 ,30874 ,11752 ,23857 ,15804 ,14728 ,22511 ,30067 ,3535 ,14993 ,27008 ,25207 ,25601 ,22739 ,15486 ,11659 ,12713 ,31106 ,10040 ,31742 ,18437 ,14800 ,20796 ,10590 ,27195 ,28679 ,13554 ,30812 ,3036 ,16032 ,5431 ,4747 ,16862 ,31234 ,18360 ,29370 ,31367 ,24920 ,20005 ,21105 ,19152 ,26353 ,8484 ,20583 ,6464 ,21422 ,4466 ,18278 ,7879 ,1448 ,4419 ,5665 ,22464 ,19792 ,12180 ,14872 ,4913 ,30788 ,31703 ,22958 ,27553 ,13616 ,25320 ,15674 ,23398 ,26043 ,5712 ,22642 ,4922 ,30102 ,9629 ,8644 ,22811 ,14139 ,6952 ,20420 ,26439 ,14866 ,5126 ,3363 ,8318 ,9067 ,16540 ,4574 ,14204 ,24085 ,24473 ,548 ,10478 ,2054 ,
      10187 ,10688 ,23757 ,25829 ,19771 ,18814 ,24295 ,17335 ,20630 ,9924 ,7506 ,3570 ,15079 ,1635 ,1777 ,5336 ,13688 ,29748 ,23793 ,31913 ,15884 ,4296 ,9228 ,21766 ,4595 ,31861 ,14349 ,20127 ,32506 ,5132 ,13607 ,22440 ,27803 ,24364 ,31444 ,30174 ,32627 ,3246 ,18854 ,21980 ,3944 ,3286 ,7079 ,18570 ,21315 ,11002 ,11415 ,4503 ,5875 ,1164 ,12052 ,13920 ,8531 ,23266 ,23495 ,12390 ,24197 ,8089 ,17420 ,25435 ,28115 ,3737 ,21632 ,31296 ,10949 ,14015 ,23907 ,19305 ,24686 ,24157 ,23724 ,7046 ,25568 ,17859 ,27520 ,31334 ,6511 ,5513 ,1352 ,12831 ,24623 ,11286 ,24719 ,12117 ,7413 ,1004 ,27140 ,24007 ,20499 ,28765 ,28717 ,24316 ,26655 ,3369 ,31694 ,30764 ,16732 ,22325 ,6261 ,27218 ,11869 ,12350 ,683 ,19646 ,25964 ,30625 ,28889 ,13135 ,21655 ,18647 ,12508 ,22065 ,21469 ,3745 ,1964 ,15714 ,10598 ,7323 ,14938 ,7724 ,16435 ,10033 ,24190 ,16924 ,4787 ,164 ,20300 ,2540 ,1495 ,32212 ,15464 ,8509 ,2802 ,14309 ,6977 ,27343 ,29892 ,19864 ,19338 ,17718 ,27033 ,9419 ,26261 ,17264 ,7131 ,6397 ,30458 ,10268 ,29000 ,4188 ,4364 ,6643 ,9751 ,6742 ,32096 ,17356 ,8857 ,8324 ,15665 ,8460 ,21212 ,7156 ,23940 ,32249 ,5925 ,4256 ,6104 ,26776 ,6361 ,20547 ,14662 ,15028 ,13297 ,25063 ,2685 ,22254 ,5900 ,18150 ,396 ,27699 ,26143 ,13713 ,29315 ,4809 ,16931 ,31977 ,21494 ,16652 ,7926 ,1956 ,30602 ,24648 ,28062 ,12841 ,22075 ,28264 ,4513 ,19731 ,10529 ,5346 ,22264 ,19244 ,3185 ,17274 ,11349 ,17213 ,25002 ,17203 ,15003 ,28813 ,27986 ,6028 ,27766 ,26363 ,14149 ,584 ,16561 ,29657 ,14048 ,10818 ,16104 ,9073 ,23389 ,18254 ,6182 ,9830 ,25714 ,27423 ,28469 ,3530 ,19147 ,22806 ,1772 ,11410 ,1347 ,12503 ,26256 ,2680 ,24997 ,24992 ,2660 ,9399 ,10982 ,5493 ,11119 ,2120 ,30047 ,21085 ,18325 ,17029 ,29857 ,3909 ,21930 ,31184 ,7814 ,15594 ,
      15579 ,21915 ,17014 ,29842 ,5478 ,2645 ,2105 ,30032 ,22791 ,28454 ,9815 ,25699 ,12488 ,1757 ,2665 ,24982 ,17188 ,11334 ,19229 ,3170 ,28249 ,28047 ,19716 ,10514 ,569 ,27751 ,28798 ,27971 ,10803 ,16546 ,9058 ,23374 ,8445 ,8842 ,6727 ,32081 ,10253 ,7116 ,4173 ,4349 ,27328 ,2787 ,32197 ,15449 ,17703 ,29877 ,9404 ,26246 ,22239 ,13282 ,20532 ,14647 ,32234 ,21197 ,4241 ,6089 ,4794 ,26128 ,18135 ,381 ,16637 ,16916 ,1941 ,30587 ,31281 ,28100 ,8074 ,17405 ,13905 ,5860 ,23251 ,23480 ,21965 ,32612 ,24349 ,31429 ,18555 ,3929 ,10987 ,11400 ,5321 ,15064 ,9909 ,7491 ,25814 ,10172 ,18799 ,24280 ,21751 ,15869 ,29733 ,23778 ,20112 ,4580 ,5117 ,13592 ,30749 ,26640 ,28750 ,28702 ,12102 ,24608 ,989 ,27125 ,7031 ,24671 ,14000 ,23892 ,31319 ,25553 ,5498 ,1337 ,22050 ,21640 ,30610 ,28874 ,27203 ,16717 ,12335 ,668 ,7709 ,10583 ,3730 ,1949 ,16909 ,16420 ,149 ,20285 ,8183 ,359 ,14778 ,25413 ,23164 ,30418 ,2159 ,29432 ,21850 ,13752 ,12974 ,19506 ,3083 ,17049 ,11124 ,27413 ,29632 ,11492 ,26688 ,30959 ,24818 ,5268 ,10894 ,23305 ,7362 ,24767 ,1547 ,25850 ,18922 ,14210 ,20411 ,9605 ,19113 ,29281 ,23690 ,9194 ,2213 ,8284 ,2577 ,31510 ,10123 ,8235 ,9526 ,22175 ,4139 ,12301 ,2125 ,6172 ,16079 ,26551 ,20987 ,32145 ,2460 ,11698 ,11231 ,20322 ,171 ,19009 ,3402 ,13488 ,26846 ,16427 ,7701 ,645 ,28664 ,20781 ,31727 ,18422 ,22724 ,26993 ,11644 ,12698 ,30859 ,2315 ,16210 ,11787 ,14713 ,11737 ,30052 ,3520 ,6003 ,6821 ,10724 ,21236 ,1127 ,19439 ,6206 ,17634 ,24494 ,27827 ,22876 ,779 ,16756 ,24091 ,26430 ,22618 ,30773 ,12165 ,5650 ,22449 ,21407 ,8469 ,18263 ,7864 ,31219 ,5416 ,30797 ,3021 ,24905 ,18345 ,21090 ,19137 ,14124 ,9614 ,22627 ,4907 ,13601 ,31688 ,15659 ,23383 ,9052 ,5111 ,20405 ,26424 ,24070 ,16525 ,533 ,10463 ,
      10448 ,24055 ,5096 ,20390 ,4892 ,14109 ,31673 ,15644 ,7849 ,21392 ,12150 ,5635 ,3006 ,31204 ,18330 ,21075 ,3505 ,14698 ,2300 ,16195 ,18407 ,28649 ,26978 ,11629 ,17619 ,1112 ,6806 ,10709 ,764 ,24479 ,24076 ,26415 ,9590 ,18907 ,24752 ,1532 ,30944 ,29617 ,5253 ,10879 ,29417 ,23149 ,344 ,14763 ,19491 ,21835 ,17034 ,11109 ,6157 ,4124 ,8220 ,9511 ,9179 ,19098 ,8269 ,2562 ,20307 ,2445 ,26536 ,20972 ,13473 ,156 ,16412 ,7686 ,30572 ,16622 ,26113 ,18120 ,14632 ,22224 ,21182 ,4226 ,4334 ,10238 ,8827 ,6712 ,15434 ,27313 ,29862 ,9389 ,24967 ,12473 ,28439 ,9800 ,29827 ,15564 ,2630 ,2090 ,10499 ,28234 ,11319 ,19214 ,27956 ,554 ,16531 ,9043 ,13577 ,20097 ,15854 ,29718 ,7476 ,5306 ,10157 ,18784 ,23465 ,13890 ,28085 ,8059 ,31414 ,21950 ,3914 ,10972 ,1322 ,31304 ,24656 ,13985 ,28687 ,30734 ,24593 ,974 ,653 ,27188 ,21625 ,30595 ,1934 ,7694 ,16405 ,134 ,119 ,1919 ,27173 ,21610 ,13970 ,1307 ,30719 ,24578 ,18769 ,7461 ,20082 ,15839 ,8044 ,23450 ,21935 ,3899 ,9374 ,15419 ,10223 ,8812 ,18105 ,30557 ,22209 ,21167 ,2075 ,29812 ,12458 ,28424 ,19199 ,10484 ,539 ,16516 ,26400 ,749 ,1097 ,6791 ,16180 ,3490 ,28634 ,26963 ,15629 ,4877 ,24040 ,5081 ,5620 ,7834 ,31189 ,18315 ,11094 ,19476 ,23134 ,329 ,1517 ,9575 ,29602 ,5238 ,2547 ,9164 ,4109 ,8205 ,20957 ,20292 ,141 ,16397 ,16382 ,20942 ,9149 ,4094 ,314 ,11079 ,9560 ,29587 ,26948 ,16165 ,734 ,1082 ,5066 ,15614 ,7819 ,31174 ,3884 ,8029 ,7446 ,20067 ,21595 ,104 ,1292 ,30704 ,21152 ,18090 ,15404 ,10208 ,28409 ,2060 ,10469 ,524 ,509 ,28394 ,18075 ,15389 ,20052 ,3869 ,89 ,1277 ,29572 ,299 ,20927 ,9134 ,1067 ,26933 ,15599 ,7804 ,7789 ,1052 ,284 ,20912 ,15374 ,494 ,3854 ,74 ,59 ,15359 ,1037 ,269 ,254 ,44 ,29 ,14 ,
      32766 ,239 ,15344 ,1022 ,20897 ,7774 ,479 ,3839 ,1262 ,20037 ,28379 ,18060 ,9119 ,29557 ,26918 ,15584 ,31159 ,5051 ,16150 ,719 ,4079 ,16367 ,11064 ,9545 ,30689 ,21580 ,8014 ,7431 ,10193 ,21137 ,2045 ,10454 ,16501 ,19184 ,29797 ,12443 ,8797 ,9359 ,30542 ,22194 ,24563 ,13955 ,1904 ,27158 ,15824 ,18754 ,23435 ,21920 ,18300 ,5605 ,4862 ,24025 ,6776 ,26385 ,3475 ,28619 ,5223 ,1502 ,19461 ,23119 ,8190 ,2532 ,20277 ,126 ,7671 ,13458 ,2430 ,26521 ,9496 ,6142 ,19083 ,8254 ,10864 ,30929 ,18892 ,24737 ,14748 ,29402 ,21820 ,17019 ,21060 ,2991 ,21377 ,12135 ,20375 ,10433 ,14094 ,31658 ,11614 ,18392 ,14683 ,2285 ,10694 ,17604 ,24464 ,24061 ,9028 ,27941 ,28219 ,11304 ,9785 ,24952 ,15549 ,2615 ,4211 ,14617 ,16607 ,26098 ,6697 ,4319 ,27298 ,29847 ,10957 ,31399 ,13875 ,28070 ,29703 ,13562 ,5291 ,10142 ,959 ,28672 ,31289 ,24641 ,30580 ,638 ,7679 ,16390 ,20270 ,16894 ,10568 ,3715 ,28859 ,22035 ,16702 ,12320 ,27110 ,12087 ,26625 ,28735 ,23877 ,7016 ,25538 ,5483 ,11385 ,18540 ,32597 ,24334 ,17390 ,31266 ,5845 ,23236 ,24265 ,25799 ,15049 ,9894 ,23763 ,21736 ,4565 ,5102 ,23359 ,10788 ,27736 ,28783 ,3155 ,17173 ,28032 ,19701 ,30017 ,5463 ,21900 ,16999 ,25684 ,22776 ,1742 ,2650 ,26231 ,17688 ,2772 ,32182 ,32066 ,8430 ,7101 ,4158 ,6074 ,32219 ,13267 ,20517 ,366 ,4779 ,16901 ,1926 ,630 ,26831 ,18994 ,3387 ,32130 ,16064 ,11683 ,11216 ,31495 ,2198 ,29266 ,23675 ,22160 ,10108 ,12286 ,2110 ,27398 ,3068 ,13737 ,12959 ,25398 ,8168 ,30403 ,2144 ,23290 ,24803 ,11477 ,26673 ,25835 ,7347 ,14195 ,20396 ,22603 ,16741 ,27812 ,22861 ,21221 ,5988 ,19424 ,6191 ,12683 ,22709 ,20766 ,31712 ,11772 ,30844 ,11722 ,30037 ,19122 ,24890 ,5401 ,30782 ,22434 ,30758 ,8454 ,18248 ,23368 ,13586 ,9599 ,22612 ,26409 ,9037 ,16510 ,518 ,
      2039 ,24458 ,4559 ,14189 ,14851 ,6937 ,3348 ,8303 ,26028 ,25305 ,22943 ,27538 ,30087 ,5697 ,8629 ,22796 ,26338 ,19990 ,29355 ,31352 ,16017 ,13539 ,4732 ,16847 ,1433 ,4451 ,20568 ,6449 ,19777 ,4404 ,14857 ,4898 ,5392 ,9268 ,30352 ,17877 ,8891 ,19824 ,28181 ,6548 ,11544 ,4664 ,13245 ,25170 ,15206 ,2927 ,23535 ,28459 ,14978 ,22496 ,23842 ,15789 ,2855 ,12659 ,18592 ,2232 ,31091 ,15471 ,25192 ,25586 ,14785 ,10025 ,10575 ,27180 ,951 ,15270 ,4006 ,5531 ,10382 ,9711 ,22121 ,31584 ,29487 ,12212 ,13802 ,8963 ,15752 ,29943 ,13385 ,9820 ,18229 ,11197 ,23217 ,19682 ,28600 ,3820 ,31639 ,2596 ,28310 ,31565 ,16828 ,6529 ,18820 ,14904 ,6943 ,14115 ,24881 ,4945 ,13047 ,17524 ,12887 ,6603 ,21544 ,31529 ,20207 ,1199 ,12753 ,1370 ,22531 ,29157 ,28912 ,25704 ,14023 ,17968 ,878 ,12849 ,8358 ,30820 ,12776 ,28329 ,15278 ,20789 ,28108 ,7919 ,16630 ,26839 ,13466 ,20950 ,2525 ,4772 ,10018 ,24175 ,15699 ,21454 ,7308 ,14923 ,19631 ,11854 ,22310 ,6246 ,13120 ,25949 ,18632 ,12493 ,12816 ,6496 ,17844 ,27505 ,19290 ,10934 ,24142 ,23709 ,23992 ,7398 ,11271 ,24704 ,24301 ,20484 ,3354 ,31679 ,22425 ,32491 ,31846 ,14334 ,31898 ,13673 ,4281 ,9213 ,17320 ,19756 ,10673 ,23742 ,3555 ,20615 ,1620 ,1762 ,4488 ,21300 ,3271 ,7064 ,30159 ,27788 ,3231 ,18839 ,12375 ,8516 ,1149 ,12037 ,25420 ,24182 ,3722 ,21617 ,24633 ,7911 ,31962 ,21479 ,27684 ,5885 ,13698 ,29300 ,26761 ,5910 ,7141 ,23925 ,15013 ,6346 ,25048 ,2670 ,17249 ,27018 ,19849 ,19323 ,8494 ,1480 ,14294 ,6962 ,6628 ,28985 ,6382 ,30443 ,17341 ,9736 ,8309 ,15650 ,18239 ,16089 ,29642 ,14033 ,6013 ,14988 ,26348 ,14134 ,5331 ,4498 ,12826 ,22060 ,17259 ,22249 ,17198 ,24987 ,24977 ,26241 ,11395 ,1332 ,27408 ,6167 ,3515 ,19132 ,21070 ,11104 ,9384 ,10967 ,3894 ,18310 ,31169 ,7799 ,
      26913 ,23430 ,21815 ,27293 ,25533 ,1737 ,12281 ,11717 ,8624 ,23530 ,13380 ,28907 ,18627 ,1615 ,25043 ,17193 ,25038 ,25487 ,7587 ,13153 ,10302 ,26075 ,25265 ,13821 ,29088 ,32454 ,25084 ,14435 ,20636 ,30231 ,26034 ,7855 ,19415 ,8751 ,433 ,30643 ,2384 ,10648 ,7633 ,8982 ,29220 ,25352 ,8408 ,12637 ,2726 ,25638 ,25492 ,11339 ,6336 ,27638 ,26302 ,21024 ,31800 ,25374 ,3308 ,2479 ,13199 ,2809 ,4686 ,25982 ,23171 ,15706 ,28866 ,13977 ,13867 ,870 ,32681 ,18665 ,30492 ,13648 ,27071 ,12231 ,3627 ,15117 ,1818 ,20700 ,30315 ,7219 ,7592 ,19234 ,26751 ,27585 ,16283 ,11923 ,11456 ,7993 ,16807 ,11250 ,6874 ,25886 ,16304 ,21673 ,9930 ,32370 ,25311 ,21398 ,5979 ,30125 ,10348 ,15983 ,3121 ,22400 ,20863 ,20341 ,12549 ,14551 ,20184 ,12526 ,2350 ,22990 ,13158 ,3175 ,23915 ,28523 ,32689 ,22083 ,23024 ,3044 ,1393 ,29506 ,4014 ,31735 ,8082 ,31970 ,26121 ,19002 ,2438 ,9157 ,5216 ,6067 ,31084 ,12368 ,13192 ,12012 ,25760 ,29962 ,17123 ,9661 ,19556 ,11962 ,30277 ,19915 ,10307 ,28254 ,31952 ,15965 ,20682 ,11905 ,14417 ,27275 ,12619 ,21006 ,27469 ,12923 ,11944 ,11887 ,7512 ,8676 ,22949 ,12156 ,22594 ,22843 ,23657 ,12941 ,9876 ,3697 ,16981 ,32164 ,23101 ,12425 ,18042 ,701 ,2267 ,26503 ,26080 ,28052 ,7901 ,17506 ,8945 ,19664 ,6431 ,14171 ,25152 ,15771 ,12019 ,14316 ,6228 ,27487 ,30425 ,21461 ,22042 ,1314 ,31391 ,17960 ,28515 ,8694 ,18488 ,21275 ,5806 ,26570 ,14481 ,14516 ,30998 ,6279 ,30894 ,22674 ,25270 ,19721 ,27674 ,19362 ,1842 ,27236 ,3209 ,3453 ,25130 ,13404 ,31022 ,5744 ,13318 ,7530 ,3576 ,19580 ,27544 ,5641 ,22852 ,22334 ,24373 ,22343 ,7165 ,30134 ,8760 ,9839 ,16234 ,23608 ,29134 ,22967 ,17795 ,12998 ,13826 ,10519 ,29290 ,4954 ,9277 ,12174 ,32500 ,26649 ,8851 ,16098 ,10797 ,20106 ,18916 ,16750 ,758 ,27950 ,19193 ,28403 ,
      21131 ,17598 ,21730 ,7341 ,4398 ,14898 ,20478 ,9730 ,30225 ,32364 ,8670 ,19574 ,32332 ,32306 ,29093 ,574 ,14284 ,26471 ,15933 ,11980 ,23576 ,27918 ,17928 ,3421 ,32422 ,1583 ,27606 ,10616 ,15085 ,32338 ,30093 ,3012 ,20757 ,29125 ,11165 ,9679 ,4632 ,9993 ,24426 ,13507 ,28953 ,6314 ,26209 ,14956 ,11822 ,20452 ,32459 ,27756 ,1470 ,18722 ,5019 ,7742 ,14585 ,606 ,13426 ,10401 ,25767 ,6984 ,17656 ,17141 ,2166 ,7315 ,16709 ,30726 ,29695 ,8350 ,23016 ,19933 ,9445 ,25924 ,32027 ,19028 ,7245 ,8566 ,5782 ,1982 ,2890 ,32396 ,25089 ,28803 ,17239 ,13100 ,15186 ,15732 ,6677 ,9099 ,25664 ,22140 ,17775 ,30257 ,2706 ,30295 ,1641 ,32312 ,5703 ,31210 ,22700 ,23599 ,27865 ,3763 ,12583 ,19606 ,11028 ,31603 ,29023 ,5158 ,13024 ,10325 ,1661 ,15907 ,14440 ,27976 ,19313 ,8702 ,18673 ,28272 ,19941 ,16040 ,24841 ,190 ,5539 ,18430 ,17413 ,21487 ,18128 ,3395 ,26529 ,4102 ,23112 ,20510 ,25579 ,12030 ,25975 ,27480 ,17134 ,16446 ,3955 ,31033 ,14492 ,24208 ,16245 ,4606 ,20641 ,10808 ,6372 ,6885 ,3638 ,16942 ,12560 ,9762 ,29903 ,4025 ,29231 ,16572 ,22275 ,13210 ,1783 ,29099 ,8635 ,18336 ,11763 ,17786 ,7256 ,10051 ,29034 ,24117 ,2953 ,5550 ,28964 ,4430 ,18371 ,25778 ,5723 ,32433 ,30236 ,16551 ,28975 ,14236 ,29183 ,29980 ,17075 ,29242 ,3966 ,26865 ,29969 ,27350 ,11566 ,16453 ,29439 ,14930 ,12327 ,24585 ,10134 ,28321 ,29498 ,182 ,20218 ,7373 ,21861 ,15289 ,11555 ,24505 ,30870 ,31102 ,31230 ,1444 ,26039 ,9063 ,17331 ,21762 ,21976 ,12386 ,7042 ,24003 ,19642 ,7720 ,27339 ,6639 ,26772 ,4805 ,5342 ,580 ,22802 ,21081 ,30028 ,10510 ,4345 ,6085 ,23476 ,24276 ,27121 ,664 ,29428 ,23301 ,31506 ,20318 ,12694 ,17630 ,7860 ,23379 ,15640 ,11625 ,10875 ,2558 ,4222 ,2086 ,18780 ,970 ,24574 ,21163 ,26959 ,5234 ,29583 ,30700 ,1273 ,70 ,
      475 ,11060 ,30538 ,3471 ,19079 ,14090 ,15545 ,5287 ,16698 ,5841 ,28028 ,7097 ,11679 ,30399 ,19420 ,8450 ,3344 ,4728 ,28177 ,18588 ,22117 ,31635 ,21540 ,12772 ,7304 ,24138 ,4277 ,3227 ,13694 ,14290 ,26344 ,3511 ,12277 ,25261 ,7629 ,3304 ,27067 ,16803 ,20859 ,1389 ,25756 ,12615 ,16977 ,25148 ,5802 ,25126 ,8756 ,8847 ,20474 ,17924 ,24422 ,13422 ,32023 ,25660 ,11024 ,24837 ,17130 ,29899 ,2949 ,3962 ,21857 ,19638 ,27117 ,18776 ,15541 ,21536 ,20855 ,11020 ,32723 ,3795 ,32727 ,1218 ,5008 ,9315 ,18018 ,1860 ,2002 ,23075 ,438 ,6732 ,23982 ,27897 ,7972 ,27254 ,8147 ,16346 ,3799 ,10913 ,18711 ,17560 ,16325 ,21333 ,29754 ,26477 ,19996 ,14704 ,10099 ,22665 ,5181 ,19380 ,916 ,18204 ,32731 ,23324 ,14574 ,8124 ,28577 ,11433 ,15506 ,23631 ,30648 ,32086 ,24694 ,18496 ,30500 ,4521 ,9453 ,5439 ,1222 ,20226 ,10390 ,22732 ,13913 ,27692 ,14640 ,32138 ,9504 ,322 ,4855 ,2765 ,23835 ,3264 ,26295 ,8938 ,5012 ,29176 ,24415 ,1693 ,3673 ,13336 ,8586 ,14391 ,2389 ,10258 ,17834 ,826 ,32555 ,7548 ,15163 ,21354 ,9319 ,26707 ,9982 ,18958 ,21694 ,32645 ,23799 ,15939 ,29361 ,2306 ,31486 ,14472 ,26189 ,5762 ,20164 ,13360 ,18022 ,30978 ,20746 ,26605 ,1884 ,18872 ,12733 ,22923 ,10653 ,7121 ,6486 ,17462 ,1700 ,21998 ,28557 ,28008 ,1864 ,22550 ,9668 ,19871 ,10746 ,31040 ,13759 ,11861 ,12094 ,7468 ,24944 ,6595 ,22392 ,19598 ,18196 ,15245 ,2006 ,11511 ,26198 ,24232 ,22570 ,31462 ,31126 ,5190 ,7638 ,4178 ,19280 ,17742 ,20724 ,30192 ,17298 ,24541 ,23079 ,28931 ,6303 ,29055 ,5946 ,3594 ,31919 ,11986 ,31358 ,16201 ,23666 ,6270 ,31453 ,24382 ,23949 ,10357 ,442 ,25723 ,11811 ,27874 ,11174 ,27562 ,7265 ,19530 ,8987 ,4354 ,23699 ,13056 ,30361 ,5659 ,31855 ,28759 ,6736 ,29651 ,27745 ,15863 ,24761 ,27821 ,1106 ,28228 ,29806 ,18084 ,
      30683 ,11608 ,24259 ,23284 ,1427 ,28304 ,23986 ,6622 ,29082 ,6868 ,27463 ,31016 ,32416 ,17769 ,29225 ,27333 ,7298 ,18705 ,9976 ,6297 ,32289 ,17581 ,27901 ,1566 ,32295 ,13083 ,25907 ,8549 ,15890 ,23582 ,16023 ,18413 ,18985 ,28506 ,22383 ,14534 ,7202 ,853 ,7976 ,25869 ,30214 ,25470 ,1720 ,23513 ,25621 ,8734 ,25357 ,2792 ,21444 ,17489 ,3680 ,12408 ,19898 ,6050 ,27258 ,12906 ,19563 ,19345 ,21258 ,14499 ,12981 ,22317 ,26632 ,20089 ,9020 ,24873 ,5971 ,22692 ,10091 ,26814 ,8151 ,24786 ,21719 ,18523 ,22018 ,12070 ,22759 ,10771 ,8413 ,32202 ,2515 ,5588 ,9342 ,13938 ,29540 ,222 ,16350 ,21563 ,17587 ,2974 ,6125 ,30912 ,4302 ,27924 ,13545 ,28655 ,26822 ,17951 ,6586 ,1182 ,29926 ,15253 ,3803 ,31548 ,4387 ,19973 ,6920 ,25288 ,2910 ,9251 ,12642 ,15454 ,24165 ,21283 ,13656 ,19739 ,25932 ,4755 ,10917 ,7381 ,9719 ,27001 ,5868 ,5893 ,22232 ,16072 ,6150 ,11087 ,5598 ,17681 ,22489 ,21293 ,27631 ,17499 ,18715 ,14229 ,17917 ,17455 ,17482 ,17438 ,25227 ,18462 ,2731 ,17708 ,22300 ,17472 ,836 ,25453 ,17752 ,11591 ,17564 ,13066 ,27907 ,5571 ,26797 ,18506 ,9234 ,17934 ,4738 ,26984 ,32121 ,18479 ,18187 ,8107 ,23058 ,21519 ,16329 ,17543 ,14273 ,4711 ,14073 ,5824 ,25109 ,25244 ,25643 ,29882 ,11844 ,17445 ,13343 ,26588 ,14374 ,2748 ,21337 ,18941 ,11969 ,17725 ,15228 ,24215 ,19513 ,6253 ,28742 ,15846 ,11296 ,17516 ,15975 ,3755 ,19372 ,1174 ,29758 ,4964 ,27595 ,18160 ,6407 ,28533 ,28823 ,27648 ,25497 ,9409 ,13110 ,25217 ,22901 ,8712 ,20593 ,18732 ,26481 ,20430 ,1572 ,14246 ,6895 ,28133 ,21772 ,3427 ,16853 ,11635 ,11207 ,26561 ,11502 ,17978 ,6831 ,22506 ,20000 ,9624 ,15074 ,21310 ,6506 ,21650 ,27028 ,13292 ,11344 ,26251 ,12483 ,17698 ,18550 ,31314 ,3078 ,4134 ,14708 ,24900 ,3001 ,19486 ,15429 ,31409 ,8039 ,5615 ,5061 ,1062 ,
      29552 ,18749 ,29397 ,4314 ,7011 ,22771 ,10103 ,30839 ,5692 ,2922 ,29938 ,29152 ,25944 ,20610 ,6341 ,22244 ,1610 ,25633 ,7214 ,22985 ,19910 ,26498 ,22669 ,12993 ,32301 ,20447 ,32391 ,15902 ,4601 ,32428 ,1439 ,17625 ,30394 ,25121 ,23070 ,23626 ,14386 ,22918 ,5185 ,19525 ,17764 ,8729 ,10766 ,9246 ,18457 ,25239 ,27643 ,13287 ,20605 ,25234 ,8593 ,21784 ,31769 ,28835 ,19384 ,8377 ,30284 ,27040 ,6843 ,16252 ,3090 ,13127 ,23884 ,8051 ,16599 ,12745 ,20176 ,13016 ,28569 ,6912 ,920 ,13771 ,15175 ,28150 ,31060 ,23811 ,14820 ,8598 ,26307 ,20537 ,17310 ,14263 ,26730 ,31931 ,27377 ,31138 ,18208 ,12795 ,13089 ,7277 ,23961 ,17813 ,31867 ,1589 ,4457 ,1118 ,8159 ,3444 ,24532 ,29766 ,4048 ,2014 ,32735 ,28348 ,6666 ,15518 ,928 ,13844 ,9465 ,21789 ,21029 ,14652 ,23732 ,5814 ,27079 ,10537 ,32035 ,16870 ,23328 ,21869 ,22129 ,11652 ,23259 ,13706 ,21190 ,11691 ,19091 ,9568 ,6769 ,32059 ,2848 ,30152 ,31793 ,6424 ,14578 ,17068 ,32016 ,28550 ,19891 ,14367 ,31762 ,31774 ,31805 ,32239 ,31836 ,18177 ,15144 ,20145 ,32004 ,19060 ,8128 ,897 ,25913 ,10072 ,32270 ,7183 ,14355 ,27612 ,20574 ,6812 ,27389 ,27665 ,19271 ,31879 ,2836 ,14832 ,28581 ,12868 ,29684 ,9477 ,4060 ,8778 ,32047 ,28840 ,25379 ,21202 ,32481 ,18469 ,14398 ,9857 ,31781 ,25514 ,11437 ,3102 ,19922 ,9426 ,23557 ,4613 ,17056 ,25956 ,7023 ,23457 ,14609 ,1191 ,14543 ,5150 ,8116 ,19965 ,15510 ,17987 ,5771 ,20828 ,17099 ,24391 ,19048 ,19389 ,3313 ,4246 ,31888 ,23048 ,26167 ,22361 ,31824 ,29775 ,23635 ,11143 ,8555 ,4981 ,9951 ,32524 ,20133 ,10622 ,6455 ,10715 ,12950 ,27227 ,30183 ,22352 ,32258 ,15992 ,30652 ,27432 ,2879 ,3772 ,9688 ,13625 ,10060 ,8382 ,2484 ,6094 ,9203 ,17533 ,17886 ,22458 ,14343 ,28711 ,32090 ,14042 ,28792 ,29727 ,1541 ,22870 ,6800 ,11313 ,12452 ,15398 ,
      7425 ,2279 ,9888 ,26667 ,6443 ,6523 ,24698 ,30437 ,14429 ,21667 ,11881 ,7524 ,10610 ,30289 ,13204 ,4799 ,3221 ,21327 ,32639 ,3588 ,8543 ,30906 ,18500 ,28127 ,15896 ,17807 ,7177 ,32518 ,32512 ,15091 ,19783 ,770 ,11468 ,13309 ,5937 ,9942 ,26155 ,30327 ,30504 ,7938 ,29012 ,2362 ,3133 ,8869 ,23036 ,27045 ,2814 ,26133 ,27778 ,2738 ,2396 ,16116 ,31812 ,11361 ,4525 ,23183 ,10314 ,26268 ,28481 ,20648 ,11131 ,18639 ,25545 ,21942 ,6689 ,22523 ,2342 ,1653 ,15498 ,2902 ,9457 ,20808 ,27854 ,1673 ,12595 ,9295 ,19953 ,6848 ,4691 ,18140 ,4478 ,11834 ,4644 ,12192 ,14597 ,20017 ,5443 ,2178 ,23588 ,9641 ,25332 ,15097 ,5138 ,32344 ,4410 ,24485 ,24794 ,5735 ,29046 ,4972 ,17087 ,11519 ,1226 ,29451 ,12572 ,17995 ,13779 ,1795 ,20816 ,16257 ,25987 ,386 ,7054 ,26578 ,12239 ,5354 ,19036 ,31242 ,20230 ,15297 ,31592 ,12706 ,23488 ,29308 ,4234 ,11224 ,8262 ,29595 ,28612 ,4151 ,2225 ,18832 ,2472 ,15764 ,10394 ,26858 ,24830 ,22543 ,12899 ,18934 ,8370 ,3095 ,23176 ,16642 ,1139 ,15218 ,8903 ,16768 ,2867 ,14725 ,22736 ,14797 ,16029 ,24917 ,21419 ,19789 ,13613 ,30099 ,14863 ,24082 ,25826 ,3567 ,31910 ,20124 ,30171 ,18567 ,13917 ,25432 ,19302 ,31331 ,12114 ,24313 ,27215 ,13132 ,15711 ,16921 ,8506 ,17715 ,10265 ,17353 ,32246 ,15025 ,27696 ,16649 ,28261 ,17271 ,6025 ,10815 ,27420 ,12500 ,5490 ,3906 ,29839 ,25696 ,3167 ,27968 ,32078 ,15446 ,14644 ,378 ,17402 ,31426 ,7488 ,23775 ,28699 ,23889 ,28871 ,1946 ,25410 ,19503 ,30956 ,25847 ,9191 ,22172 ,32142 ,13485 ,18419 ,11784 ,21233 ,776 ,22446 ,3018 ,4904 ,26421 ,20387 ,5632 ,16192 ,10706 ,1529 ,14760 ,9508 ,20969 ,18117 ,6709 ,9797 ,19211 ,29715 ,8056 ,13982 ,30592 ,21607 ,15836 ,8809 ,28421 ,6788 ,5078 ,326 ,8202 ,4091 ,1079 ,20064 ,10205 ,15386 ,9131 ,20909 ,266 ,
      15341 ,28376 ,16147 ,8011 ,29794 ,1901 ,4859 ,19458 ,2427 ,18889 ,21374 ,14680 ,28216 ,16604 ,13872 ,31286 ,10565 ,26622 ,32594 ,15046 ,27733 ,21897 ,2769 ,13264 ,18991 ,29263 ,13734 ,11474 ,27809 ,20763 ,5398 ,9596 ,4556 ,22940 ,29352 ,20565 ,30349 ,13242 ,23839 ,25189 ,4003 ,13799 ,23214 ,16825 ,13044 ,12750 ,875 ,28105 ,10015 ,22307 ,17841 ,11268 ,31843 ,10670 ,3268 ,1146 ,31959 ,7138 ,19846 ,6379 ,29639 ,12823 ,11392 ,9381 ,21812 ,13377 ,7584 ,25081 ,430 ,8405 ,26299 ,4683 ,32678 ,1815 ,16280 ,16301 ,10345 ,20181 ,32686 ,8079 ,31081 ,19553 ,20679 ,11941 ,23654 ,18039 ,8942 ,6225 ,28512 ,30995 ,1839 ,13315 ,24370 ,29131 ,9274 ,18913 ,21727 ,8667 ,15930 ,27603 ,11162 ,26206 ,5016 ,17653 ,23013 ,5779 ,15183 ,2703 ,27862 ,13021 ,18670 ,17410 ,25576 ,14489 ,3635 ,22272 ,7253 ,18368 ,29180 ,11563 ,29495 ,30867 ,21973 ,26769 ,4342 ,31503 ,10872 ,26956 ,30535 ,28025 ,28174 ,4274 ,7626 ,16974 ,24419 ,2946 ,20852 ,18015 ,7969 ,16322 ,5178 ,28574 ,30497 ,13910 ,23832 ,3670 ,32552 ,21691 ,26186 ,1881 ,1697 ,10743 ,22389 ,22567 ,20721 ,5943 ,31450 ,11171 ,30358 ,24758 ,24256 ,27460 ,9973 ,25904 ,22380 ,1717 ,3677 ,21255 ,5968 ,22015 ,9339 ,6122 ,6583 ,6917 ,13653 ,5865 ,22486 ,17479 ,833 ,26794 ,18184 ,14070 ,13340 ,15225 ,15972 ,6404 ,22898 ,6892 ,11499 ,6503 ,18547 ,15426 ,29394 ,29935 ,7211 ,32388 ,23067 ,10763 ,8590 ,6840 ,20173 ,31057 ,26727 ,23958 ,24529 ,925 ,27076 ,23256 ,2845 ,19888 ,15141 ,32267 ,19268 ,4057 ,14395 ,23554 ,14540 ,17096 ,26164 ,9948 ,30180 ,9685 ,17883 ,1538 ,9885 ,11878 ,32636 ,7174 ,5934 ,3130 ,2393 ,28478 ,2339 ,12592 ,4641 ,25329 ,29043 ,13776 ,12236 ,23485 ,2222 ,12896 ,8900 ,21416 ,31907 ,12111 ,10262 ,6022 ,3164 ,7485 ,30953 ,21230 ,16189 ,9794 ,8806 ,20061 ,
      16144 ,21371 ,32591 ,13731 ,29349 ,23211 ,17838 ,19843 ,7581 ,16277 ,20676 ,1836 ,15927 ,15180 ,3632 ,21970 ,28171 ,7966 ,32549 ,20718 ,9970 ,9336 ,830 ,22895 ,7208 ,26724 ,15138 ,26161 ,32633 ,4638 ,8897 ,30950 ,32588 ,20673 ,32546 ,15135 ,32543 ,32572 ,32559 ,798 ,3616 ,7565 ,32575 ,29333 ,814 ,28155 ,15122 ,32617 ,19814 ,843 ,32562 ,4827 ,15151 ,10840 ,7552 ,8910 ,20689 ,30465 ,801 ,3645 ,26695 ,17851 ,32604 ,10230 ,10856 ,29479 ,3619 ,7237 ,5000 ,21711 ,15167 ,27846 ,32670 ,32662 ,7568 ,414 ,8926 ,31065 ,1823 ,24354 ,5382 ,18975 ,32578 ,27717 ,4843 ,15325 ,21358 ,28200 ,859 ,3987 ,29336 ,30333 ,3252 ,9999 ,19830 ,29623 ,18531 ,15956 ,817 ,18168 ,3661 ,24240 ,9323 ,6567 ,30481 ,20836 ,28158 ,7610 ,1681 ,23816 ,20705 ,31434 ,17867 ,14524 ,15125 ,19252 ,8574 ,29378 ,26711 ,24513 ,12220 ,2323 ,32620 ,5918 ,10246 ,2206 ,30937 ,16173 ,9352 ,17166 ,19817 ,13666 ,10641 ,3690 ,9986 ,24110 ,16796 ,13353 ,846 ,21512 ,22911 ,14825 ,30320 ,18560 ,13235 ,1710 ,32565 ,16670 ,20734 ,16478 ,18962 ,30371 ,7982 ,26886 ,4830 ,30510 ,18860 ,24432 ,28187 ,5259 ,17381 ,14408 ,15154 ,31995 ,26177 ,16677 ,21698 ,17896 ,26740 ,26007 ,10843 ,27089 ,14460 ,8603 ,7224 ,3934 ,4654 ,25460 ,7555 ,12249 ,20152 ,2406 ,32649 ,16775 ,11912 ,10275 ,8913 ,16949 ,30966 ,27512 ,24341 ,8819 ,24729 ,8955 ,20692 ,1974 ,1852 ,12062 ,23803 ,9287 ,16293 ,406 ,30468 ,32699 ,27996 ,26312 ,7597 ,10992 ,15196 ,25611 ,804 ,18683 ,6474 ,5029 ,15943 ,26449 ,25875 ,29193 ,3648 ,7944 ,21986 ,13513 ,6554 ,10885 ,23227 ,20997 ,26698 ,888 ,10734 ,23852 ,29365 ,22637 ,9919 ,3281 ,17854 ,30620 ,19859 ,20542 ,19239 ,11405 ,28449 ,2782 ,32607 ,24666 ,13747 ,8230 ,2310 ,5411 ,21387 ,23144 ,10233 ,13885 ,7456 ,4872 ,16160 ,294 ,
      1257 ,24558 ,10859 ,4206 ,27105 ,30012 ,31490 ,12678 ,26023 ,11539 ,29482 ,20202 ,19626 ,17315 ,26756 ,5326 ,8619 ,29215 ,3622 ,12544 ,17118 ,23096 ,14476 ,16229 ,30220 ,28948 ,7240 ,29018 ,3950 ,28959 ,11550 ,29423 ,16693 ,25751 ,5003 ,14569 ,24410 ,20741 ,26193 ,11806 ,29077 ,30209 ,21714 ,4382 ,17912 ,14268 ,27590 ,15069 ,5687 ,17759 ,15170 ,6661 ,32011 ,29679 ,5766 ,2874 ,14424 ,29007 ,27849 ,12567 ,24825 ,19297 ,17397 ,18112 ,2422 ,3998 ,32673 ,23008 ,20847 ,5963 ,20168 ,2334 ,7576 ,3611 ,32665 ,30476 ,16791 ,26735 ,16288 ,9914 ,26018 ,29072 ,7571 ,10286 ,12265 ,26897 ,13364 ,18611 ,25476 ,29204 ,417 ,2368 ,3292 ,6320 ,4670 ,23155 ,22026 ,12003 ,8929 ,6415 ,16965 ,22578 ,18026 ,2251 ,10291 ,17107 ,31068 ,13176 ,12603 ,31936 ,11928 ,7496 ,27528 ,31006 ,1826 ,3193 ,5790 ,31375 ,30982 ,30878 ,13810 ,16218 ,24357 ,7149 ,8835 ,29274 ,18900 ,742 ,16494 ,23352 ,5385 ,22418 ,19408 ,22587 ,20750 ,11756 ,12270 ,31479 ,18978 ,32114 ,30387 ,27382 ,11461 ,25819 ,4549 ,24249 ,32581 ,17374 ,16686 ,20254 ,26609 ,23861 ,1726 ,30001 ,27720 ,3139 ,7085 ,26215 ,13251 ,350 ,20261 ,5207 ,4846 ,6760 ,30526 ,16485 ,1888 ,15808 ,26902 ,1246 ,15328 ,20881 ,11048 ,31143 ,7998 ,10177 ,24448 ,11598 ,21361 ,20359 ,19067 ,7655 ,18876 ,14732 ,27282 ,4195 ,28203 ,9769 ,5275 ,10941 ,31273 ,30564 ,13450 ,15262 ,862 ,8342 ,21528 ,24865 ,12737 ,22515 ,13369 ,29471 ,3990 ,10366 ,31623 ,18213 ,16812 ,18804 ,14841 ,1417 ,29339 ,16001 ,3332 ,2023 ,22927 ,30071 ,23519 ,11528 ,30336 ,8875 ,18576 ,14962 ,25176 ,14769 ,3706 ,12359 ,3255 ,30143 ,4265 ,22409 ,10657 ,3539 ,18616 ,19615 ,10002 ,15683 ,24126 ,12800 ,11255 ,24285 ,8293 ,6612 ,19833 ,8478 ,13682 ,24617 ,7125 ,14997 ,17182 ,5315 ,29626 ,5997 ,3499 ,24961 ,9368 ,3878 ,
      5045 ,2985 ,18534 ,3062 ,19984 ,11191 ,6490 ,27012 ,25481 ,27579 ,15959 ,19356 ,26465 ,13094 ,6879 ,21756 ,4722 ,27891 ,820 ,17736 ,18699 ,5582 ,17466 ,25211 ,25627 ,14257 ,18171 ,23042 ,21321 ,11828 ,15212 ,19497 ,26616 ,19547 ,3664 ,19882 ,7960 ,18969 ,1704 ,25605 ,29209 ,29066 ,24243 ,1411 ,27885 ,7282 ,25891 ,15874 ,13529 ,17571 ,9326 ,29524 ,8135 ,9004 ,22002 ,22743 ,12626 ,4371 ,6570 ,29910 ,10901 ,24149 ,5852 ,22216 ,9488 ,10374 ,30484 ,9437 ,32715 ,10083 ,28561 ,15490 ,422 ,4992 ,20839 ,32707 ,3783 ,23966 ,16309 ,29738 ,26328 ,7288 ,28161 ,22101 ,15529 ,459 ,28012 ,11663 ,8740 ,25740 ,7613 ,27051 ,11008 ,20458 ,2933 ,21841 ,12078 ,9652 ,1684 ,28541 ,18006 ,31470 ,1868 ,12717 ,2373 ,24399 ,23819 ,26279 ,9303 ,17818 ,21678 ,23783 ,31342 ,6287 ,20708 ,17282 ,1990 ,24928 ,22554 ,31110 ,8971 ,11795 ,31437 ,23933 ,6720 ,23683 ,24745 ,1090 ,12436 ,28776 ,17870 ,14327 ,30636 ,12934 ,9672 ,10044 ,3297 ,5755 ,14527 ,8100 ,23619 ,31872 ,9935 ,20117 ,20558 ,25897 ,15128 ,31988 ,14562 ,6753 ,19875 ,31746 ,25363 ,29668 ,19255 ,2820 ,11421 ,32465 ,23541 ,17040 ,23868 ,30268 ,8577 ,31753 ,5169 ,30378 ,10750 ,18441 ,6325 ,5676 ,29381 ,6995 ,22653 ,1594 ,32375 ,4585 ,4441 ,13073 ,26714 ,27361 ,904 ,16583 ,31044 ,14804 ,21013 ,6650 ,24516 ,4032 ,23312 ,23716 ,23243 ,21174 ,8246 ,31576 ,12223 ,19020 ,1210 ,24778 ,13763 ,20800 ,4675 ,27838 ,2326 ,15482 ,5427 ,4462 ,25316 ,5122 ,19767 ,15880 ,32623 ,8527 ,24682 ,7409 ,11865 ,10594 ,2798 ,28996 ,5921 ,26139 ,4509 ,27762 ,28465 ,11115 ,5474 ,28245 ,10249 ,32230 ,13901 ,25810 ,12098 ,27199 ,23160 ,24814 ,2209 ,2456 ,22720 ,1123 ,21403 ,13597 ,4888 ,18403 ,30940 ,9175 ,14628 ,29823 ,7472 ,28683 ,13966 ,18101 ,16176 ,1513 ,310 ,21591 ,20048 ,15370 ,
      7770 ,16363 ,9355 ,26381 ,6138 ,10429 ,24948 ,13558 ,22031 ,31262 ,17169 ,8426 ,16060 ,8164 ,5984 ,30754 ,6933 ,13535 ,19820 ,12655 ,9707 ,3816 ,6599 ,30816 ,21450 ,10930 ,13669 ,27784 ,5881 ,1476 ,14984 ,6163 ,1733 ,26071 ,10644 ,25370 ,13644 ,7989 ,22396 ,3040 ,12008 ,27271 ,3693 ,14167 ,21271 ,3449 ,30130 ,26645 ,14894 ,27914 ,9989 ,602 ,25920 ,9095 ,19602 ,16036 ,27476 ,9758 ,24113 ,29238 ,7369 ,23999 ,24272 ,2082 ,14086 ,31631 ,16799 ,25656 ,3791 ,16342 ,18200 ,5435 ,8934 ,21350 ,13356 ,28004 ,15241 ,24537 ,10353 ,28755 ,28300 ,17577 ,849 ,6046 ,26810 ,218 ,15249 ,4751 ,17495 ,11587 ,21515 ,2744 ,1170 ,18728 ,22502 ,4130 ,22767 ,26494 ,22914 ,28831 ,6908 ,31134 ,2010 ,16866 ,6420 ,19056 ,14828 ,25510 ,19961 ,29771 ,15988 ,28707 ,6519 ,30902 ,30323 ,11357 ,2898 ,20013 ,11515 ,31238 ,15760 ,14721 ,18563 ,15021 ,15442 ,22168 ,14756 ,5074 ,1897 ,21893 ,13238 ,10666 ,8401 ,18035 ,26202 ,18364 ,16970 ,1877 ,1713 ,14066 ,10759 ,4053 ,3126 ,12107 ,23207 ,9332 ,32568 ,10836 ,21707 ,15321 ,24236 ,29374 ,3686 ,16474 ,16673 ,2402 ,12058 ,5025 ,23848 ,8226 ,30008 ,23092 ,20737 ,29675 ,5959 ,26893 ,22574 ,31371 ,22583 ,20250 ,16481 ,7651 ,24861 ,2019 ,22405 ,24613 ,11187 ,5578 ,18965 ,9000 ,10079 ,455 ,31466 ,24924 ,12930 ,6749 ,30374 ,16579 ,24774 ,7405 ,25806 ,29819 ,10425 ,3812 ,7985 ,9091 ,16338 ,214 ,31130 ,20009 ,18031 ,15317 ,26889 ,451 ,210 ,32740 ,20868 ,994 ,28590 ,29530 ,4833 ,30661 ,2503 ,32744 ,5194 ,21109 ,12414 ,1235 ,30513 ,16122 ,13926 ,7748 ,15795 ,9517 ,16990 ,692 ,18863 ,8769 ,6113 ,20872 ,7642 ,19156 ,2256 ,11037 ,24435 ,23407 ,2962 ,28353 ,20346 ,27130 ,2586 ,21553 ,28190 ,18272 ,4290 ,998 ,4182 ,26357 ,28041 ,10166 ,5262 ,19433 ,28643 ,15558 ,30551 ,98 ,
      4073 ,20369 ,17384 ,25392 ,16011 ,28594 ,19284 ,8488 ,10296 ,11450 ,14411 ,3203 ,23570 ,6671 ,12554 ,7036 ,22111 ,8141 ,15157 ,17292 ,32283 ,29534 ,17746 ,20587 ,19904 ,27371 ,31998 ,31818 ,8537 ,14591 ,2861 ,9185 ,27727 ,23648 ,26180 ,19262 ,9964 ,4837 ,20728 ,6468 ,17112 ,12259 ,16680 ,3326 ,18693 ,15523 ,14556 ,24676 ,9701 ,26804 ,21701 ,2497 ,32277 ,30665 ,30196 ,21426 ,11951 ,32103 ,17899 ,22282 ,1554 ,11278 ,15056 ,12465 ,21052 ,18221 ,26743 ,17231 ,23974 ,2507 ,17302 ,4470 ,31073 ,5374 ,26010 ,26320 ,28292 ,933 ,20189 ,14005 ,941 ,9010 ,10846 ,21042 ,30671 ,32748 ,24545 ,18282 ,6056 ,23341 ,27092 ,11367 ,23272 ,612 ,12665 ,19104 ,10779 ,22834 ,14463 ,27656 ,27451 ,5198 ,23083 ,7883 ,13181 ,19397 ,8606 ,25020 ,6856 ,13849 ,12531 ,23897 ,5521 ,22682 ,7227 ,17221 ,32404 ,21113 ,28935 ,1452 ,29951 ,11745 ,3937 ,6354 ,27321 ,10116 ,29410 ,15622 ,13948 ,5456 ,4657 ,19749 ,25345 ,12418 ,6307 ,4423 ,12608 ,26598 ,25463 ,4704 ,8722 ,9470 ,2355 ,31324 ,13792 ,22008 ,7558 ,26000 ,30202 ,1239 ,29059 ,5669 ,27264 ,20243 ,12252 ,4531 ,23501 ,13432 ,18598 ,8275 ,3146 ,9867 ,20155 ,2827 ,22371 ,30517 ,5950 ,22468 ,31941 ,4538 ,2409 ,10547 ,28494 ,21794 ,22995 ,25558 ,12202 ,18513 ,32652 ,5364 ,7190 ,16126 ,3598 ,19796 ,11894 ,17363 ,16778 ,13217 ,25857 ,24711 ,9901 ,28431 ,12127 ,19674 ,11915 ,15724 ,27246 ,13930 ,31923 ,12184 ,11933 ,27709 ,10278 ,22093 ,6038 ,21034 ,13163 ,5503 ,15742 ,22749 ,8916 ,28282 ,21432 ,7752 ,11990 ,14876 ,12912 ,29990 ,16952 ,23189 ,12396 ,10407 ,2238 ,2568 ,19692 ,32155 ,30969 ,12859 ,21246 ,15799 ,31362 ,4917 ,7501 ,7074 ,27515 ,28884 ,19333 ,14657 ,3180 ,1342 ,9810 ,32192 ,24344 ,13995 ,12969 ,9521 ,16205 ,30792 ,12145 ,339 ,8822 ,28080 ,20077 ,24035 ,729 ,20922 ,
      18055 ,27153 ,24732 ,26093 ,28730 ,16994 ,23670 ,31707 ,27533 ,25165 ,8958 ,1365 ,6241 ,23737 ,23920 ,22055 ,28902 ,12632 ,20695 ,12521 ,11957 ,696 ,6274 ,22962 ,19569 ,14951 ,1977 ,10320 ,24203 ,25773 ,31097 ,20313 ,7092 ,25143 ,1855 ,11428 ,13331 ,18867 ,31457 ,27557 ,31011 ,23508 ,12065 ,25283 ,17433 ,5819 ,28528 ,21645 ,29147 ,9241 ,23806 ,13839 ,14362 ,8773 ,24386 ,13620 ,7519 ,8864 ,9290 ,1790 ,18929 ,24308 ,23770 ,19206 ,14675 ,16820 ,16296 ,2698 ,16317 ,6117 ,23953 ,25324 ,1831 ,29328 ,409 ,7605 ,21507 ,27084 ,32694 ,30615 ,20197 ,4377 ,30471 ,13171 ,32109 ,20876 ,10361 ,15678 ,19351 ,1406 ,32702 ,26274 ,8095 ,6990 ,15477 ,2451 ,8421 ,14162 ,27999 ,25505 ,14061 ,7646 ,446 ,23402 ,3198 ,3321 ,26315 ,25015 ,4699 ,10542 ,22088 ,28879 ,1360 ,25278 ,7600 ,25010 ,25097 ,19160 ,25727 ,26047 ,13393 ,30060 ,10995 ,25056 ,29870 ,12294 ,21828 ,7827 ,15817 ,25677 ,15199 ,3548 ,2719 ,2260 ,11815 ,5716 ,5795 ,12726 ,25614 ,25102 ,18450 ,32040 ,23029 ,27208 ,13037 ,6576 ,807 ,14453 ,17905 ,11041 ,27878 ,22646 ,21264 ,24854 ,18686 ,28487 ,17426 ,17662 ,25198 ,26542 ,26222 ,7892 ,6477 ,32472 ,22477 ,24439 ,11178 ,4926 ,31380 ,13439 ,5032 ,19165 ,17669 ,16875 ,3049 ,16722 ,4935 ,17941 ,15946 ,22824 ,27619 ,23411 ,27566 ,30106 ,8683 ,8331 ,26452 ,29106 ,14217 ,20491 ,21743 ,10491 ,18384 ,31557 ,25878 ,30249 ,17552 ,2966 ,7269 ,9633 ,30987 ,3979 ,29196 ,25732 ,11579 ,23333 ,1398 ,12340 ,12877 ,29916 ,3651 ,27441 ,22288 ,28357 ,19534 ,8648 ,14505 ,29460 ,7947 ,20654 ,25441 ,17147 ,25592 ,20978 ,32173 ,19655 ,21989 ,9848 ,26785 ,20350 ,8991 ,22815 ,30883 ,31612 ,13516 ,26052 ,5559 ,21874 ,29511 ,673 ,31519 ,31538 ,6557 ,7873 ,9222 ,27134 ,4358 ,14143 ,19710 ,18793 ,10888 ,6200 ,26972 ,2624 ,22203 ,1286 ,
      9539 ,31652 ,23230 ,2138 ,16841 ,2590 ,23703 ,6956 ,13815 ,11244 ,21000 ,13398 ,3415 ,22134 ,4019 ,7714 ,12766 ,10907 ,26701 ,28925 ,1560 ,21557 ,13060 ,20424 ,12987 ,12789 ,891 ,11137 ,28121 ,2172 ,14791 ,13479 ,13258 ,6219 ,10737 ,23548 ,22889 ,28194 ,30365 ,26443 ,16223 ,18605 ,23855 ,30065 ,25205 ,11657 ,31740 ,10588 ,30810 ,4745 ,29368 ,21103 ,20581 ,18276 ,5663 ,14870 ,22956 ,15672 ,22640 ,8642 ,20418 ,3361 ,4572 ,546 ,10686 ,18812 ,9922 ,1633 ,29746 ,4294 ,31859 ,5130 ,24362 ,3244 ,3284 ,11000 ,1162 ,23264 ,8087 ,3735 ,14013 ,24155 ,17857 ,5511 ,11284 ,1002 ,28763 ,3367 ,22323 ,12348 ,30623 ,18645 ,3743 ,7321 ,10031 ,162 ,32210 ,14307 ,19862 ,9417 ,6395 ,4186 ,6740 ,8322 ,7154 ,4254 ,20545 ,25061 ,18148 ,13711 ,31975 ,1954 ,12839 ,19729 ,19242 ,17211 ,28811 ,26361 ,29655 ,9071 ,9828 ,3528 ,11408 ,2678 ,9397 ,2118 ,17027 ,31182 ,21913 ,2643 ,28452 ,1755 ,11332 ,28045 ,27749 ,16544 ,8840 ,7114 ,2785 ,29875 ,13280 ,21195 ,26126 ,16914 ,28098 ,5858 ,32610 ,3927 ,15062 ,10170 ,15867 ,4578 ,26638 ,24606 ,24669 ,25551 ,21638 ,16715 ,10581 ,16418 ,357 ,30416 ,13750 ,17047 ,11490 ,5266 ,24765 ,14208 ,29279 ,8282 ,8233 ,12299 ,26549 ,11696 ,19007 ,16425 ,20779 ,26991 ,2313 ,11735 ,6819 ,19437 ,27825 ,24089 ,12163 ,8467 ,5414 ,18343 ,9612 ,31686 ,5109 ,16523 ,24053 ,14107 ,21390 ,31202 ,14696 ,28647 ,1110 ,24477 ,18905 ,29615 ,23147 ,21833 ,4122 ,19096 ,2443 ,154 ,16620 ,22222 ,10236 ,27311 ,12471 ,15562 ,28232 ,552 ,20095 ,5304 ,13888 ,21948 ,31302 ,30732 ,27186 ,7692 ,1917 ,1305 ,7459 ,23448 ,15417 ,30555 ,29810 ,10482 ,747 ,3488 ,4875 ,7832 ,19474 ,9573 ,9162 ,20290 ,20940 ,11077 ,16163 ,15612 ,8027 ,102 ,18088 ,2058 ,28392 ,3867 ,297 ,26931 ,1050 ,492 ,15357 ,42 ,
      32764 ,20895 ,1260 ,9117 ,31157 ,4077 ,30687 ,10191 ,16499 ,8795 ,24561 ,15822 ,18298 ,6774 ,5221 ,8188 ,7669 ,9494 ,10862 ,14746 ,21058 ,20373 ,11612 ,10692 ,9026 ,9783 ,4209 ,6695 ,10955 ,29701 ,957 ,30578 ,20268 ,28857 ,27108 ,23875 ,11383 ,17388 ,24263 ,23761 ,23357 ,3153 ,30015 ,25682 ,26229 ,32064 ,6072 ,364 ,628 ,32128 ,31493 ,22158 ,27396 ,25396 ,23288 ,25833 ,22601 ,21219 ,12681 ,11770 ,19120 ,22432 ,23366 ,26407 ,2037 ,14849 ,26026 ,30085 ,26336 ,16015 ,1431 ,19775 ,5390 ,8889 ,11542 ,15204 ,14976 ,2853 ,31089 ,14783 ,949 ,10380 ,29485 ,15750 ,18227 ,28598 ,28308 ,18818 ,24879 ,12885 ,20205 ,22529 ,14021 ,8356 ,15276 ,16628 ,2523 ,15697 ,19629 ,13118 ,12814 ,19288 ,23990 ,24299 ,22423 ,31896 ,17318 ,3553 ,4486 ,30157 ,12373 ,25418 ,24631 ,27682 ,26759 ,15011 ,17247 ,8492 ,6626 ,17339 ,18237 ,6011 ,5329 ,17257 ,24975 ,27406 ,21068 ,3892 ,26911 ,25531 ,8622 ,18625 ,25036 ,10300 ,29086 ,20634 ,19413 ,2382 ,29218 ,2724 ,6334 ,31798 ,13197 ,23169 ,13865 ,30490 ,3625 ,30313 ,26749 ,11454 ,6872 ,9928 ,5977 ,3119 ,12547 ,2348 ,23913 ,23022 ,4012 ,26119 ,5214 ,13190 ,17121 ,30275 ,31950 ,14415 ,27467 ,7510 ,22592 ,9874 ,23099 ,2265 ,7899 ,6429 ,12017 ,30423 ,31389 ,18486 ,14479 ,30892 ,27672 ,3207 ,31020 ,3574 ,22850 ,7163 ,16232 ,17793 ,29288 ,32498 ,10795 ,756 ,21129 ,4396 ,30223 ,32330 ,14282 ,23574 ,32420 ,15083 ,20755 ,4630 ,28951 ,11820 ,1468 ,14583 ,25765 ,2164 ,29693 ,9443 ,7243 ,2888 ,17237 ,6675 ,17773 ,1639 ,22698 ,12581 ,29021 ,1659 ,19311 ,19939 ,5537 ,18126 ,23110 ,25973 ,3953 ,16243 ,6370 ,12558 ,29229 ,1781 ,11761 ,29032 ,28962 ,5721 ,28973 ,17073 ,29967 ,29437 ,10132 ,20216 ,11553 ,31228 ,17329 ,7040 ,27337 ,5340 ,30026 ,23474 ,29426 ,12692 ,15638 ,4220 ,24572 ,29581 ,
      473 ,19077 ,16696 ,11677 ,3342 ,22115 ,7302 ,13692 ,12275 ,27065 ,25754 ,5800 ,20472 ,32021 ,17128 ,21855 ,15539 ,32721 ,5006 ,2000 ,23980 ,8145 ,18709 ,29752 ,10097 ,914 ,14572 ,15504 ,24692 ,9451 ,10388 ,14638 ,4853 ,26293 ,24413 ,8584 ,17832 ,15161 ,9980 ,23797 ,31484 ,20162 ,20744 ,12731 ,6484 ,28555 ,9666 ,13757 ,24942 ,18194 ,26196 ,31124 ,19278 ,17296 ,6301 ,31917 ,23664 ,23947 ,11809 ,7263 ,23697 ,31853 ,27743 ,1104 ,30681 ,1425 ,29080 ,32414 ,7296 ,32287 ,32293 ,15888 ,18983 ,7200 ,30212 ,25619 ,21442 ,19896 ,19561 ,12979 ,9018 ,10089 ,21717 ,22757 ,2513 ,29538 ,17585 ,4300 ,26820 ,29924 ,4385 ,2908 ,24163 ,25930 ,9717 ,22230 ,5596 ,27629 ,17915 ,25225 ,22298 ,17750 ,27905 ,9232 ,32119 ,23056 ,14271 ,25107 ,11842 ,14372 ,11967 ,19511 ,11294 ,19370 ,27593 ,28821 ,13108 ,20591 ,1570 ,21770 ,11205 ,6829 ,15072 ,27026 ,12481 ,3076 ,2999 ,8037 ,29550 ,7009 ,5690 ,25942 ,1608 ,19908 ,32299 ,4599 ,30392 ,14384 ,17762 ,18455 ,20603 ,31767 ,30282 ,3088 ,16597 ,28567 ,15173 ,14818 ,17308 ,27375 ,13087 ,31865 ,8157 ,4046 ,6664 ,9463 ,23730 ,32033 ,22127 ,21188 ,6767 ,31791 ,32014 ,31760 ,31834 ,32002 ,25911 ,14353 ,27387 ,2834 ,29682 ,32045 ,32479 ,31779 ,19920 ,17054 ,14607 ,8114 ,5769 ,19046 ,31886 ,31822 ,8553 ,20131 ,12948 ,32256 ,2877 ,10058 ,9201 ,14341 ,28790 ,6798 ,7423 ,6441 ,14427 ,10608 ,3219 ,8541 ,15894 ,32510 ,11466 ,26153 ,29010 ,23034 ,27776 ,31810 ,10312 ,11129 ,6687 ,15496 ,27852 ,19951 ,4476 ,14595 ,23586 ,5136 ,24792 ,17085 ,12570 ,20814 ,7052 ,19034 ,31590 ,4232 ,28610 ,2470 ,24828 ,8368 ,1137 ,2865 ,16027 ,13611 ,25824 ,30169 ,19300 ,27213 ,8504 ,32244 ,28259 ,27418 ,29837 ,32076 ,17400 ,28697 ,25408 ,9189 ,18417 ,22444 ,20385 ,1527 ,18115 ,29713 ,21605 ,6786 ,4089 ,15384 ,
      15339 ,29792 ,2425 ,28214 ,10563 ,27731 ,18989 ,27807 ,4554 ,30347 ,4001 ,13042 ,10013 ,31841 ,31957 ,29637 ,21810 ,428 ,32676 ,10343 ,31079 ,23652 ,28510 ,24368 ,21725 ,11160 ,23011 ,27860 ,25574 ,7251 ,29493 ,4340 ,30533 ,7624 ,20850 ,5176 ,23830 ,26184 ,22387 ,31448 ,24254 ,22378 ,5966 ,6581 ,22484 ,18182 ,15970 ,11497 ,29392 ,23065 ,20171 ,24527 ,2843 ,19266 ,14538 ,30178 ,9883 ,5932 ,2337 ,29041 ,2220 ,31905 ,3162 ,16187 ,16142 ,29347 ,7579 ,15925 ,28169 ,9968 ,7206 ,32631 ,32586 ,32541 ,3614 ,812 ,19812 ,15149 ,20687 ,26693 ,10854 ,4998 ,32668 ,8924 ,5380 ,4841 ,857 ,3250 ,18529 ,3659 ,30479 ,1679 ,17865 ,8572 ,12218 ,10244 ,9350 ,10639 ,16794 ,22909 ,13233 ,20732 ,7980 ,18858 ,17379 ,26175 ,26738 ,14458 ,4652 ,20150 ,11910 ,30964 ,24727 ,1850 ,16291 ,27994 ,15194 ,6472 ,25873 ,21984 ,23225 ,10732 ,9917 ,19857 ,28447 ,13745 ,21385 ,7454 ,1255 ,27103 ,26021 ,19624 ,8617 ,17116 ,30218 ,3948 ,16691 ,24408 ,29075 ,17910 ,5685 ,32009 ,14422 ,24823 ,2420 ,20845 ,7574 ,16789 ,26016 ,12263 ,25474 ,3290 ,22024 ,16963 ,10289 ,12601 ,27526 ,5788 ,13808 ,8833 ,16492 ,19406 ,12268 ,30385 ,4547 ,16684 ,1724 ,7083 ,20259 ,30524 ,26900 ,11046 ,24446 ,19065 ,27280 ,5273 ,13448 ,21526 ,13367 ,31621 ,14839 ,3330 ,23517 ,18574 ,3704 ,4263 ,18614 ,24124 ,8291 ,13680 ,17180 ,3497 ,5043 ,19982 ,25479 ,26463 ,4720 ,18697 ,25625 ,21319 ,26614 ,7958 ,29207 ,27883 ,13527 ,8133 ,12624 ,10899 ,9486 ,32713 ,420 ,3781 ,26326 ,15527 ,8738 ,11006 ,12076 ,18004 ,2371 ,9301 ,31340 ,1988 ,8969 ,6718 ,12434 ,30634 ,3295 ,23617 ,20556 ,14560 ,25361 ,11419 ,23866 ,5167 ,6323 ,22651 ,4439 ,902 ,21011 ,23310 ,8244 ,1208 ,4673 ,5425 ,19765 ,24680 ,2796 ,4507 ,5472 ,13899 ,23158 ,22718 ,4886 ,14626 ,13964 ,308 ,
      7768 ,6136 ,22029 ,16058 ,6931 ,9705 ,21448 ,5879 ,1731 ,13642 ,12006 ,21269 ,14892 ,25918 ,27474 ,7367 ,14084 ,3789 ,8932 ,15239 ,28298 ,26808 ,17493 ,1168 ,22765 ,6906 ,6418 ,19959 ,6517 ,2896 ,15758 ,15440 ,1895 ,8399 ,16968 ,10757 ,23205 ,21705 ,3684 ,12056 ,30006 ,5957 ,22581 ,24859 ,11185 ,10077 ,12928 ,24772 ,10423 ,16336 ,18029 ,208 ,28588 ,2501 ,12412 ,13924 ,16988 ,6111 ,2254 ,2960 ,2584 ,4288 ,28039 ,28641 ,4071 ,16009 ,10294 ,23568 ,22109 ,32281 ,19902 ,8535 ,27725 ,9962 ,17110 ,18691 ,9699 ,32275 ,11949 ,1552 ,21050 ,23972 ,31071 ,28290 ,939 ,30669 ,6054 ,23270 ,10777 ,27449 ,13179 ,6854 ,5519 ,32402 ,29949 ,27319 ,13946 ,25343 ,12606 ,8720 ,13790 ,30200 ,27262 ,23499 ,3144 ,22369 ,31939 ,28492 ,12200 ,7188 ,11892 ,25855 ,12125 ,27244 ,11931 ,6036 ,15740 ,21430 ,12910 ,12394 ,19690 ,21244 ,7499 ,19331 ,9808 ,12967 ,12143 ,20075 ,18053 ,28728 ,27531 ,6239 ,28900 ,11955 ,19567 ,24201 ,7090 ,13329 ,31009 ,17431 ,29145 ,14360 ,7517 ,18927 ,14673 ,16315 ,1829 ,21505 ,20195 ,32107 ,19349 ,8093 ,8419 ,14059 ,3196 ,4697 ,1358 ,25095 ,13391 ,29868 ,15815 ,2717 ,5793 ,18448 ,13035 ,17903 ,21262 ,17424 ,26220 ,22475 ,31378 ,17667 ,4933 ,27617 ,8681 ,14215 ,18382 ,17550 ,30985 ,11577 ,12875 ,22286 ,14503 ,25439 ,32171 ,26783 ,30881 ,5557 ,31517 ,9220 ,19708 ,26970 ,9537 ,16839 ,13813 ,3413 ,12764 ,1558 ,12985 ,28119 ,13256 ,22887 ,16221 ,25203 ,30808 ,20579 ,22954 ,20416 ,10684 ,29744 ,24360 ,1160 ,14011 ,11282 ,22321 ,3741 ,32208 ,6393 ,7152 ,18146 ,12837 ,28809 ,9826 ,9395 ,21911 ,11330 ,8838 ,13278 ,28096 ,15060 ,26636 ,21636 ,355 ,11488 ,29277 ,26547 ,20777 ,6817 ,12161 ,9610 ,24051 ,14694 ,18903 ,4120 ,16618 ,12469 ,20093 ,31300 ,1915 ,15415 ,745 ,19472 ,20938 ,8025 ,28390 ,1048 ,
      32762 ,31155 ,16497 ,18296 ,7667 ,21056 ,9024 ,10953 ,20266 ,11381 ,23355 ,26227 ,626 ,27394 ,22599 ,19118 ,2035 ,26334 ,5388 ,14974 ,947 ,18225 ,24877 ,14019 ,2521 ,12812 ,22421 ,4484 ,24629 ,17245 ,18235 ,24973 ,26909 ,25034 ,19411 ,6332 ,13863 ,26747 ,5975 ,23911 ,5212 ,31948 ,22590 ,7897 ,31387 ,27670 ,22848 ,29286 ,21127 ,14280 ,20753 ,1466 ,29691 ,17235 ,22696 ,19309 ,23108 ,6368 ,11759 ,28971 ,10130 ,17327 ,30024 ,15636 ,471 ,3340 ,12273 ,20470 ,15537 ,23978 ,10095 ,24690 ,4851 ,17830 ,31482 ,6482 ,24940 ,19276 ,23662 ,23695 ,30679 ,7294 ,18981 ,21440 ,9016 ,2511 ,26818 ,24161 ,5594 ,22296 ,32117 ,11840 ,11292 ,13106 ,11203 ,12479 ,29548 ,1606 ,30390 ,20601 ,16595 ,17306 ,8155 ,23728 ,6765 ,31832 ,27385 ,32477 ,14605 ,31884 ,12946 ,9199 ,7421 ,3217 ,11464 ,27774 ,6685 ,4474 ,24790 ,7050 ,28608 ,1135 ,25822 ,8502 ,29835 ,25406 ,20383 ,21603 ,15337 ,10561 ,4552 ,10011 ,21808 ,31077 ,21723 ,25572 ,30531 ,23828 ,24252 ,22482 ,29390 ,2841 ,9881 ,2218 ,16140 ,28167 ,32584 ,19810 ,10852 ,5378 ,18527 ,17863 ,9348 ,13231 ,17377 ,4650 ,24725 ,15192 ,23223 ,28445 ,1253 ,8615 ,16689 ,5683 ,2418 ,26014 ,22022 ,27524 ,16490 ,4545 ,20257 ,24444 ,13446 ,14837 ,3702 ,8289 ,5041 ,4718 ,26612 ,13525 ,9484 ,26324 ,12074 ,31338 ,12432 ,20554 ,23864 ,4437 ,8242 ,19763 ,5470 ,4884 ,7766 ,6929 ,1729 ,14890 ,14082 ,28296 ,22763 ,6515 ,1893 ,23203 ,30004 ,11183 ,10421 ,28586 ,16986 ,2582 ,4069 ,22107 ,27723 ,9697 ,21048 ,937 ,10775 ,5517 ,13944 ,13788 ,3142 ,12198 ,12123 ,15738 ,19688 ,9806 ,18051 ,28898 ,7088 ,29143 ,14671 ,20193 ,8417 ,1356 ,15813 ,13033 ,26218 ,4931 ,18380 ,12873 ,32169 ,31515 ,9535 ,12762 ,13254 ,30806 ,10682 ,14009 ,32206 ,12835 ,21909 ,28094 ,353 ,20775 ,24049 ,16616 ,1913 ,20936 ,
      32760 ,7665 ,20264 ,624 ,2033 ,945 ,2519 ,24627 ,26907 ,13861 ,5210 ,31385 ,21125 ,29689 ,23106 ,10128 ,469 ,15535 ,4849 ,24938 ,30677 ,9014 ,5592 ,11290 ,29546 ,16593 ,6763 ,14603 ,7419 ,6683 ,28606 ,29833 ,15335 ,21806 ,30529 ,29388 ,16138 ,10850 ,9346 ,24723 ,1251 ,2416 ,16488 ,13444 ,5039 ,9482 ,12430 ,8240 ,7764 ,14080 ,1891 ,10419 ,4067 ,21046 ,13942 ,12121 ,18049 ,14669 ,15811 ,18378 ,9533 ,10680 ,21907 ,24047 ,32758 ,2031 ,26905 ,21123 ,467 ,30675 ,29544 ,7417 ,15333 ,16136 ,1249 ,5037 ,7762 ,4065 ,18047 ,9531 ,32756 ,465 ,15331 ,7760 ,32754 ,32752 ,226 ,1008 ,228 ,28365 ,20884 ,20023 ,1010 ,9105 ,3826 ,15570 ,230 ,23421 ,11051 ,18740 ,28367 ,24549 ,16354 ,27144 ,20886 ,29783 ,31146 ,19170 ,20025 ,8783 ,706 ,22180 ,1012 ,3461 ,8001 ,26371 ,9107 ,18286 ,21567 ,24011 ,3828 ,19447 ,10180 ,1488 ,15572 ,8176 ,10441 ,112 ,232 ,16887 ,24451 ,4765 ,23423 ,6060 ,17591 ,20503 ,11053 ,2758 ,11601 ,17674 ,18742 ,32052 ,2272 ,4144 ,28369 ,28018 ,21364 ,17159 ,24551 ,23345 ,2978 ,28769 ,16356 ,21886 ,20362 ,5449 ,27146 ,25670 ,31645 ,2636 ,20888 ,25524 ,19070 ,7002 ,29785 ,27096 ,6129 ,28721 ,31148 ,10554 ,7658 ,16880 ,19172 ,28845 ,26508 ,12306 ,20027 ,5831 ,18879 ,31252 ,8785 ,11371 ,30916 ,24320 ,708 ,15035 ,14735 ,25785 ,22182 ,23749 ,17006 ,5088 ,1014 ,14181 ,27285 ,7333 ,3463 ,23276 ,4306 ,26659 ,8003 ,13723 ,4198 ,3054 ,26373 ,25384 ,26085 ,2130 ,9109 ,11669 ,28206 ,16050 ,18288 ,616 ,27928 ,3373 ,21569 ,29252 ,9772 ,2184 ,24013 ,22146 ,2602 ,2096 ,3830 ,11708 ,5278 ,30830 ,19449 ,12669 ,13549 ,31698 ,10182 ,27798 ,10944 ,16727 ,1490 ,21207 ,28057 ,6177 ,15574 ,8440 ,31276 ,30744 ,8178 ,19108 ,28659 ,30768 ,10443 ,9585 ,30567 ,13572 ,114 ,26395 ,16377 ,504 ,
      234 ,19179 ,13453 ,27936 ,16889 ,10783 ,26826 ,16736 ,24453 ,9263 ,15265 ,4940 ,4767 ,32486 ,7906 ,16084 ,23425 ,8746 ,865 ,30120 ,6062 ,22838 ,17955 ,22329 ,17593 ,29120 ,8345 ,23594 ,20505 ,17781 ,28316 ,10505 ,11055 ,25256 ,21531 ,22660 ,2760 ,14467 ,6590 ,6265 ,11603 ,28501 ,24868 ,17946 ,17676 ,18474 ,17511 ,26556 ,18744 ,25116 ,12740 ,3439 ,32054 ,27660 ,1186 ,27222 ,2274 ,13304 ,22518 ,5730 ,4146 ,3562 ,25691 ,5627 ,28371 ,22935 ,13372 ,8662 ,28020 ,27455 ,29930 ,11873 ,21366 ,20668 ,29474 ,15951 ,17161 ,14403 ,8950 ,20992 ,24553 ,25746 ,3993 ,11998 ,23347 ,5202 ,15257 ,12354 ,2980 ,19542 ,10369 ,9647 ,28771 ,30263 ,31571 ,28240 ,16358 ,26066 ,31626 ,26489 ,21888 ,23087 ,3807 ,687 ,20364 ,23643 ,18216 ,22829 ,5451 ,9862 ,19669 ,32150 ,27148 ,25138 ,16815 ,14157 ,25672 ,7887 ,31552 ,19650 ,31647 ,6214 ,18807 ,14302 ,2638 ,30411 ,14102 ,1300 ,20890 ,28852 ,14844 ,15692 ,25526 ,13185 ,4391 ,25968 ,19072 ,26288 ,1420 ,27624 ,7004 ,31786 ,6436 ,2465 ,29787 ,7619 ,29342 ,10634 ,27098 ,19401 ,19977 ,30629 ,6131 ,8394 ,16004 ,25338 ,28723 ,2712 ,16834 ,11325 ,31150 ,25029 ,3335 ,1601 ,10556 ,8610 ,6924 ,28893 ,7660 ,21801 ,2026 ,23416 ,16882 ,25519 ,14176 ,11703 ,19174 ,25251 ,22930 ,26061 ,28847 ,25024 ,25292 ,13139 ,26510 ,25070 ,30074 ,32440 ,12308 ,20622 ,22783 ,7841 ,20029 ,25297 ,23522 ,32356 ,5833 ,6860 ,2914 ,21659 ,18881 ,16269 ,11531 ,27571 ,31254 ,11442 ,25157 ,11236 ,8787 ,27057 ,30339 ,13634 ,11373 ,13853 ,9255 ,18651 ,30918 ,1804 ,8878 ,15103 ,24322 ,30301 ,6535 ,19220 ,710 ,13144 ,18579 ,22976 ,15037 ,12535 ,12646 ,12512 ,14737 ,10334 ,14965 ,30111 ,25787 ,3107 ,15776 ,20327 ,22184 ,1379 ,25179 ,3030 ,23751 ,23901 ,15458 ,22069 ,17008 ,8068 ,14772 ,31721 ,5090 ,26107 ,27167 ,9143 ,
      1016 ,26515 ,3709 ,3381 ,14183 ,5525 ,24169 ,21473 ,27287 ,18659 ,12362 ,8688 ,7335 ,19927 ,12024 ,176 ,3465 ,11014 ,3258 ,19592 ,23278 ,22686 ,21287 ,3749 ,4308 ,13010 ,30146 ,5144 ,26661 ,1647 ,18826 ,27962 ,8005 ,25075 ,4268 ,32382 ,13725 ,7231 ,13660 ,1968 ,4200 ,23002 ,22412 ,8336 ,3056 ,9431 ,14321 ,19014 ,26375 ,25650 ,10660 ,9085 ,25386 ,17225 ,19743 ,15718 ,26087 ,2692 ,3542 ,30243 ,2132 ,1627 ,1749 ,31196 ,9111 ,30079 ,18619 ,32324 ,11671 ,32408 ,25936 ,10602 ,28208 ,15919 ,19618 ,26457 ,16052 ,23562 ,6233 ,3407 ,18290 ,20464 ,10005 ,14884 ,618 ,21117 ,4759 ,7327 ,27930 ,8656 ,15686 ,32350 ,3375 ,32318 ,14910 ,560 ,21571 ,32445 ,24129 ,20438 ,29254 ,28939 ,10921 ,14942 ,9774 ,11151 ,12803 ,29111 ,2186 ,4618 ,27492 ,13493 ,24015 ,13412 ,11258 ,592 ,22148 ,1456 ,7385 ,7728 ,2604 ,17642 ,24288 ,6970 ,2098 ,2152 ,31666 ,30712 ,3832 ,12313 ,8296 ,14916 ,11710 ,29955 ,9723 ,16439 ,5280 ,29169 ,6615 ,14222 ,30832 ,17061 ,30430 ,26851 ,19451 ,2939 ,19836 ,24103 ,12671 ,11749 ,27005 ,10037 ,13551 ,18357 ,8481 ,4416 ,31700 ,5709 ,6949 ,16537 ,10184 ,20627 ,13685 ,4592 ,27800 ,3941 ,5872 ,24194 ,10946 ,25565 ,24620 ,20496 ,16729 ,25961 ,21466 ,16432 ,1492 ,29889 ,7128 ,9748 ,21209 ,6358 ,5897 ,16928 ,28059 ,22261 ,15000 ,16558 ,6179 ,1769 ,2657 ,18322 ,15576 ,22788 ,17185 ,566 ,8442 ,27325 ,22236 ,4791 ,31278 ,21962 ,5318 ,21748 ,30746 ,7028 ,22047 ,7706 ,8180 ,21847 ,29629 ,7359 ,19110 ,10120 ,16076 ,168 ,28661 ,30856 ,6000 ,24491 ,30770 ,31216 ,14121 ,9049 ,10445 ,7846 ,3502 ,17616 ,9587 ,29414 ,6154 ,20304 ,30569 ,4331 ,24964 ,10496 ,13574 ,23462 ,1319 ,650 ,116 ,18766 ,9371 ,2072 ,26397 ,15626 ,11091 ,2544 ,16379 ,26945 ,3881 ,21149 ,506 ,29569 ,7786 ,56 ,
      236 ,20034 ,5048 ,21577 ,19181 ,13952 ,5602 ,1499 ,13455 ,30926 ,2988 ,18389 ,27938 ,14614 ,31396 ,28669 ,16891 ,12084 ,18537 ,25796 ,10785 ,5460 ,17685 ,32216 ,26828 ,2195 ,3065 ,24800 ,16738 ,22706 ,24887 ,13583 ,24455 ,25302 ,19987 ,4448 ,9265 ,4661 ,22493 ,15468 ,15267 ,12209 ,11194 ,31562 ,4942 ,1196 ,17965 ,20786 ,4769 ,11851 ,6493 ,7395 ,32488 ,19753 ,21297 ,8513 ,7908 ,5907 ,27015 ,28982 ,16086 ,4495 ,26238 ,11101 ,23427 ,23527 ,25484 ,32451 ,8748 ,25349 ,27635 ,2806 ,867 ,15114 ,27582 ,25883 ,30122 ,14548 ,28520 ,31732 ,6064 ,9658 ,15962 ,12920 ,22840 ,12422 ,17503 ,14313 ,17957 ,14513 ,19359 ,5741 ,22331 ,23605 ,4951 ,20103 ,17595 ,32361 ,26468 ,1580 ,29122 ,6311 ,18719 ,6981 ,8347 ,8563 ,13097 ,30254 ,23596 ,5155 ,8699 ,18427 ,20507 ,31030 ,6882 ,16569 ,17783 ,4427 ,14233 ,27347 ,28318 ,24502 ,21759 ,6636 ,10507 ,23298 ,11622 ,21160 ,11057 ,5838 ,4725 ,24135 ,25258 ,12612 ,17921 ,29896 ,21533 ,9312 ,27894 ,17557 ,22662 ,8121 ,18493 ,22729 ,2762 ,1690 ,823 ,18955 ,14469 ,26602 ,17459 ,19868 ,6592 ,24229 ,17739 ,29052 ,6267 ,27871 ,13053 ,15860 ,11605 ,6865 ,18702 ,13080 ,28503 ,25467 ,17486 ,19342 ,24870 ,18520 ,5585 ,2971 ,17948 ,19970 ,21280 ,26998 ,17678 ,17452 ,17469 ,5568 ,18476 ,4708 ,17442 ,17722 ,17513 ,18157 ,25214 ,14243 ,26558 ,21307 ,17695 ,19483 ,18746 ,2919 ,25630 ,20444 ,25118 ,8726 ,25231 ,27037 ,12742 ,28147 ,14260 ,7274 ,3441 ,15515 ,5811 ,11649 ,32056 ,28547 ,18174 ,10069 ,27662 ,9474 ,18466 ,9423 ,1188 ,20825 ,23045 ,4978 ,27224 ,3769 ,17530 ,29724 ,2276 ,21664 ,21324 ,17804 ,13306 ,2359 ,2735 ,26265 ,22520 ,1670 ,11831 ,9638 ,5732 ,17992 ,26575 ,12703 ,4148 ,22540 ,15215 ,24914 ,3564 ,31328 ,17712 ,17268 ,25693 ,31423 ,19500 ,11781 ,5629 ,6706 ,15833 ,1076 ,
      28373 ,18886 ,26619 ,29260 ,22937 ,13796 ,22304 ,7135 ,13374 ,1812 ,19550 ,30992 ,8664 ,5776 ,14486 ,30864 ,28022 ,18012 ,3667 ,22564 ,27457 ,22012 ,17476 ,6401 ,29932 ,31054 ,19885 ,17093 ,11875 ,12589 ,12893 ,7482 ,21368 ,16274 ,7963 ,26721 ,20670 ,7562 ,840 ,30462 ,29476 ,32659 ,18972 ,3984 ,15953 ,20833 ,14521 ,2320 ,17163 ,13350 ,1707 ,26883 ,14405 ,26004 ,25457 ,10272 ,8952 ,403 ,25608 ,29190 ,20994 ,3278 ,2779 ,23141 ,24555 ,11536 ,29212 ,28945 ,25748 ,30206 ,17756 ,29004 ,3995 ,3608 ,29069 ,29201 ,12000 ,17104 ,31003 ,16215 ,23349 ,31476 ,24246 ,29998 ,5204 ,1243 ,11595 ,4192 ,15259 ,29468 ,1414 ,11525 ,12356 ,19612 ,6609 ,5312 ,2982 ,27576 ,27888 ,14254 ,19544 ,29063 ,17568 ,4368 ,10371 ,4989 ,7285 ,25737 ,9649 ,24396 ,6284 ,11792 ,28773 ,5752 ,25894 ,29665 ,30265 ,5673 ,13070 ,6647 ,31573 ,27835 ,15877 ,28993 ,28242 ,24811 ,18400 ,18098 ,16360 ,31259 ,13532 ,10927 ,26068 ,27268 ,27911 ,9755 ,31628 ,21347 ,17574 ,11584 ,26491 ,19053 ,30899 ,14718 ,21890 ,1874 ,9329 ,16471 ,23089 ,20247 ,5575 ,6746 ,3809 ,15314 ,29527 ,1232 ,689 ,11034 ,21550 ,10163 ,20366 ,11447 ,8138 ,27368 ,23645 ,12256 ,26801 ,32100 ,18218 ,5371 ,9007 ,23338 ,22831 ,19394 ,22679 ,11742 ,5453 ,26595 ,22005 ,20240 ,9864 ,4535 ,18510 ,17360 ,19671 ,27706 ,22746 ,29987 ,32152 ,7071 ,32189 ,336 ,27150 ,25162 ,12629 ,14948 ,25140 ,23505 ,9238 ,8861 ,16817 ,29325 ,4374 ,1403 ,14159 ,3318 ,25275 ,30057 ,25674 ,12723 ,6573 ,24851 ,7889 ,13436 ,17938 ,8328 ,31554 ,3976 ,29913 ,29457 ,19652 ,31609 ,31535 ,18790 ,31649 ,11241 ,10904 ,12786 ,6216 ,18602 ,4742 ,15669 ,18809 ,3241 ,24152 ,12345 ,14304 ,4251 ,19726 ,3525 ,2640 ,7111 ,5855 ,24603 ,30413 ,8279 ,26988 ,8464 ,14104 ,29612 ,22219 ,5301 ,1302 ,3485 ,11074 ,3864 ,
      20892 ,8792 ,9491 ,9780 ,28854 ,3150 ,32125 ,21216 ,14846 ,8886 ,10377 ,12882 ,15694 ,31893 ,27679 ,6008 ,25528 ,2379 ,30487 ,3116 ,13187 ,9871 ,18483 ,7160 ,4393 ,4627 ,9440 ,12578 ,25970 ,29029 ,20213 ,23471 ,19074 ,27062 ,32718 ,911 ,26290 ,20159 ,18191 ,23944 ,1422 ,7197 ,10086 ,29921 ,27626 ,23053 ,19367 ,6826 ,7006 ,14381 ,28564 ,4043 ,31788 ,2831 ,8111 ,32253 ,6438 ,26150 ,15493 ,17082 ,2467 ,30166 ,32073 ,1524 ,29789 ,30344 ,425 ,11157 ,7621 ,22375 ,23062 ,5929 ,29344 ,32538 ,4995 ,3656 ,10636 ,26172 ,1847 ,10729 ,27100 ,24405 ,20842 ,16960 ,19403 ,30521 ,21523 ,4260 ,19979 ,7955 ,32710 ,18001 ,30631 ,5164 ,1205 ,13896 ,6133 ,13639 ,3786 ,6903 ,8396 ,5954 ,16333 ,6108 ,16006 ,9959 ,23969 ,27446 ,25340 ,22366 ,27241 ,21241 ,28725 ,13326 ,16312 ,14056 ,2714 ,22472 ,17547 ,26780 ,16836 ,22884 ,29741 ,6390 ,11327 ,11485 ,14691 ,15412 ,31152 ,11378 ,26331 ,12809 ,25031 ,31945 ,14277 ,6365 ,3337 ,17827 ,7291 ,22293 ,1603 ,31829 ,3214 ,1132 ,10558 ,23825 ,28164 ,13228 ,8612 ,4542 ,4715 ,20551 ,6926 ,23200 ,22104 ,13785 ,28895 ,13030 ,12759 ,28091 ,7662 ,13858 ,15532 ,16590 ,21803 ,2413 ,14077 ,14666 ,2028 ,16133 ,462 ,28362 ,23418 ,29780 ,3458 ,19444 ,16884 ,2755 ,28015 ,21883 ,25521 ,10551 ,5828 ,15032 ,14178 ,13720 ,11666 ,29249 ,11705 ,27795 ,8437 ,9582 ,19176 ,9260 ,8743 ,29117 ,25253 ,28498 ,25113 ,13301 ,22932 ,20665 ,25743 ,19539 ,26063 ,23640 ,25135 ,6211 ,28849 ,26285 ,7616 ,8391 ,25026 ,21798 ,25248 ,25067 ,25294 ,16266 ,27054 ,1801 ,13141 ,10331 ,1376 ,8065 ,26512 ,18656 ,11011 ,13007 ,25072 ,22999 ,25647 ,2689 ,30076 ,15916 ,20461 ,8653 ,32442 ,11148 ,13409 ,17639 ,12310 ,29166 ,2936 ,18354 ,20624 ,25562 ,29886 ,22258 ,22785 ,21959 ,21844 ,30853 ,7843 ,4328 ,18763 ,26942 ,
      20031 ,30923 ,12081 ,2192 ,25299 ,12206 ,11848 ,5904 ,23524 ,15111 ,9655 ,14510 ,32358 ,8560 ,31027 ,24499 ,5835 ,9309 ,1687 ,24226 ,6862 ,18517 ,17449 ,18154 ,2916 ,28144 ,28544 ,20822 ,21661 ,1667 ,22537 ,31420 ,18883 ,1809 ,18009 ,31051 ,16271 ,32656 ,13347 ,400 ,11533 ,3605 ,31473 ,29465 ,27573 ,4986 ,5749 ,27832 ,31256 ,21344 ,1871 ,15311 ,11444 ,5368 ,26592 ,27703 ,25159 ,29322 ,12720 ,3973 ,11238 ,3238 ,7108 ,29609 ,8789 ,8883 ,2376 ,4624 ,27059 ,7194 ,14378 ,26147 ,30341 ,32535 ,24402 ,7952 ,13636 ,9956 ,13323 ,22881 ,11375 ,17824 ,23822 ,23197 ,13855 ,16130 ,2752 ,13717 ,9257 ,20662 ,26282 ,16263 ,18653 ,15913 ,29163 ,21956 ,30920 ,15108 ,9306 ,28141 ,1806 ,3602 ,21341 ,29319 ,8880 ,32532 ,17821 ,20659 ,15105 ,32529 ,7535 ,784 ,24324 ,7538 ,21681 ,10826 ,30303 ,19800 ,18945 ,4813 ,6537 ,787 ,23786 ,30451 ,19222 ,26681 ,2293 ,10216 ,712 ,24327 ,31345 ,27498 ,13146 ,11898 ,11973 ,16935 ,18581 ,7541 ,6290 ,25446 ,22978 ,20138 ,3581 ,16761 ,15039 ,21684 ,20711 ,16663 ,12537 ,17367 ,17729 ,31981 ,12648 ,10829 ,17285 ,25993 ,12514 ,14446 ,28918 ,3920 ,14739 ,30306 ,1993 ,14811 ,10336 ,16782 ,15232 ,21498 ,14967 ,19803 ,24931 ,17152 ,30113 ,10627 ,19585 ,24096 ,25789 ,18948 ,22557 ,16464 ,3109 ,13221 ,24219 ,16656 ,15778 ,4816 ,31113 ,26872 ,20329 ,18846 ,4165 ,5245 ,22186 ,6540 ,8974 ,13499 ,1381 ,25861 ,19517 ,7930 ,25181 ,790 ,11798 ,25597 ,3032 ,6460 ,27549 ,26435 ,23753 ,23789 ,31440 ,12048 ,23903 ,24715 ,6257 ,1960 ,15460 ,30454 ,23936 ,392 ,22071 ,27982 ,25710 ,10978 ,17010 ,19225 ,6723 ,20528 ,8070 ,9905 ,28746 ,30606 ,14774 ,26684 ,23686 ,20983 ,31723 ,10720 ,5646 ,22623 ,5092 ,2296 ,24748 ,8216 ,26109 ,28435 ,15850 ,24652 ,27169 ,10219 ,1093 ,23130 ,9145 ,7442 ,18071 ,280 ,
      1018 ,715 ,12439 ,24021 ,26517 ,12131 ,11300 ,28066 ,3711 ,24330 ,28779 ,32178 ,3383 ,12955 ,22857 ,30778 ,14185 ,31348 ,17873 ,15785 ,5527 ,19678 ,17520 ,12845 ,24171 ,27501 ,14330 ,7060 ,21475 ,19319 ,14029 ,1328 ,27289 ,13149 ,30639 ,21020 ,18661 ,11919 ,15979 ,22079 ,12364 ,11901 ,12937 ,19660 ,8690 ,27232 ,22339 ,12170 ,7337 ,11976 ,9675 ,7738 ,19929 ,15728 ,3759 ,28268 ,12026 ,16938 ,10047 ,29976 ,178 ,12382 ,6081 ,2554 ,3467 ,18584 ,3300 ,13418 ,11016 ,27250 ,19376 ,4517 ,3260 ,7544 ,5758 ,21994 ,19594 ,30188 ,24378 ,5655 ,23280 ,6293 ,14530 ,12404 ,22688 ,13934 ,1178 ,19735 ,21289 ,25449 ,8103 ,26584 ,3751 ,8708 ,17974 ,31310 ,4310 ,22981 ,23622 ,21780 ,13012 ,31927 ,29762 ,10533 ,30148 ,20141 ,31875 ,9853 ,5146 ,22357 ,22348 ,22454 ,26663 ,3584 ,9938 ,16112 ,1649 ,12188 ,4968 ,5350 ,18828 ,16764 ,20120 ,17349 ,27964 ,25843 ,10702 ,28417 ,8007 ,15042 ,20561 ,11264 ,25077 ,11937 ,27599 ,22268 ,4270 ,21687 ,25900 ,26790 ,32384 ,32263 ,7170 ,21412 ,13727 ,20714 ,15131 ,4823 ,7233 ,27713 ,18164 ,19248 ,13662 ,16666 ,31991 ,12245 ,1970 ,18679 ,884 ,24662 ,4202 ,12540 ,14565 ,6657 ,23004 ,10282 ,6411 ,3189 ,22414 ,17370 ,6756 ,20355 ,8338 ,15997 ,30139 ,8474 ,3058 ,17732 ,19878 ,29520 ,9433 ,22097 ,28537 ,17278 ,14323 ,31984 ,31749 ,27357 ,19016 ,8523 ,32226 ,9171 ,26377 ,12651 ,25366 ,598 ,25652 ,6042 ,28827 ,11353 ,10662 ,10832 ,29671 ,8996 ,9087 ,30657 ,8765 ,18268 ,25388 ,17288 ,19258 ,2493 ,17227 ,21038 ,27652 ,17217 ,19745 ,25996 ,2823 ,5360 ,15720 ,28278 ,12855 ,13991 ,26089 ,12517 ,11424 ,13835 ,2694 ,13167 ,25501 ,25006 ,3544 ,14449 ,32468 ,22820 ,30245 ,27437 ,9844 ,7869 ,2134 ,28921 ,23544 ,21099 ,1629 ,5507 ,9413 ,17207 ,1751 ,3923 ,17043 ,11731 ,31198 ,27307 ,23444 ,15608 ,
      9113 ,14742 ,23871 ,22154 ,30081 ,15746 ,13114 ,15007 ,18621 ,30309 ,30271 ,30888 ,32326 ,2884 ,16239 ,31224 ,11673 ,1996 ,8580 ,31120 ,32410 ,22753 ,25221 ,28817 ,25938 ,14814 ,31756 ,19042 ,10604 ,19947 ,8364 ,28693 ,28210 ,10339 ,5172 ,24523 ,15921 ,8920 ,22905 ,27990 ,19620 ,16785 ,30381 ,31617 ,26459 ,3777 ,23613 ,5421 ,16054 ,15235 ,10753 ,204 ,23564 ,28286 ,8716 ,6032 ,6235 ,21501 ,18444 ,11573 ,3409 ,1156 ,13274 ,4116 ,18292 ,14970 ,6328 ,1462 ,20466 ,21436 ,20597 ,27770 ,10007 ,19806 ,5679 ,13521 ,14886 ,9693 ,29139 ,30802 ,620 ,24934 ,29384 ,10415 ,21119 ,7756 ,18736 ,26367 ,4761 ,17155 ,6998 ,31248 ,7329 ,16046 ,30826 ,30740 ,27932 ,30116 ,22656 ,3435 ,8658 ,11994 ,26485 ,14153 ,15688 ,10630 ,1597 ,26057 ,32352 ,13630 ,22972 ,3026 ,3377 ,19588 ,32378 ,9081 ,32320 ,14880 ,20434 ,588 ,14912 ,24099 ,4588 ,9744 ,562 ,7355 ,17612 ,2068 ,21573 ,25792 ,4444 ,7391 ,32447 ,12916 ,1576 ,16565 ,24131 ,18951 ,13076 ,5564 ,20440 ,10065 ,17800 ,24910 ,29256 ,22560 ,26717 ,26879 ,28941 ,29994 ,14250 ,29661 ,10923 ,16467 ,27364 ,20236 ,14944 ,24847 ,12782 ,24599 ,9776 ,3112 ,907 ,4039 ,11153 ,16956 ,6899 ,14052 ,12805 ,13224 ,16586 ,21879 ,29113 ,8387 ,13003 ,18350 ,2188 ,24222 ,31047 ,15307 ,4620 ,23193 ,28137 ,10822 ,27494 ,16659 ,14807 ,16460 ,13495 ,12044 ,20524 ,8212 ,24017 ,15781 ,21016 ,7734 ,13414 ,12400 ,21776 ,16108 ,11260 ,4819 ,6653 ,29516 ,594 ,2489 ,13831 ,21095 ,22150 ,31116 ,24519 ,200 ,1458 ,10411 ,3431 ,9077 ,7387 ,26875 ,4035 ,15303 ,7730 ,196 ,28335 ,980 ,2606 ,20332 ,23315 ,28339 ,17644 ,2242 ,16857 ,23393 ,24290 ,18849 ,23719 ,678 ,6972 ,6099 ,10524 ,19142 ,2100 ,4168 ,23246 ,984 ,2154 ,2572 ,11639 ,18258 ,31668 ,5248 ,21177 ,10152 ,30714 ,28629 ,9555 ,84 ,
      3834 ,22189 ,8249 ,2610 ,12315 ,19696 ,11211 ,6186 ,8298 ,6543 ,31579 ,31524 ,14918 ,9208 ,29295 ,14129 ,11712 ,8977 ,12226 ,20336 ,29957 ,32159 ,26565 ,9834 ,9725 ,13502 ,19023 ,31598 ,16441 ,5545 ,15284 ,659 ,5282 ,1384 ,1213 ,23319 ,29171 ,30973 ,11506 ,25718 ,6617 ,25864 ,24781 ,31543 ,14224 ,17538 ,4959 ,9619 ,30834 ,19520 ,13766 ,28343 ,17063 ,12863 ,17982 ,27427 ,30432 ,7933 ,20803 ,29446 ,26853 ,25427 ,373 ,20964 ,19453 ,25184 ,4678 ,17648 ,2941 ,21250 ,6835 ,28473 ,19838 ,793 ,27841 ,6562 ,24105 ,17891 ,9282 ,22632 ,12673 ,11801 ,2329 ,2246 ,11751 ,15803 ,22510 ,3534 ,27007 ,25600 ,15485 ,12712 ,10039 ,18436 ,20795 ,27194 ,13553 ,3035 ,5430 ,16861 ,18359 ,31366 ,20004 ,19151 ,8483 ,6463 ,4465 ,7878 ,4418 ,22463 ,12179 ,4912 ,31702 ,27552 ,25319 ,23397 ,5711 ,4921 ,9628 ,22810 ,6951 ,26438 ,5125 ,8317 ,16539 ,14203 ,24472 ,10477 ,10186 ,23756 ,19770 ,24294 ,20629 ,7505 ,15078 ,1776 ,13687 ,23792 ,15883 ,9227 ,4594 ,14348 ,32505 ,13606 ,27802 ,31443 ,32626 ,18853 ,3943 ,7078 ,21314 ,11414 ,5874 ,12051 ,8530 ,23494 ,24196 ,17419 ,28114 ,21631 ,10948 ,23906 ,24685 ,23723 ,25567 ,27519 ,6510 ,1351 ,24622 ,24718 ,7412 ,27139 ,20498 ,28716 ,26654 ,31693 ,16731 ,6260 ,11868 ,682 ,25963 ,28888 ,21654 ,12507 ,21468 ,1963 ,10597 ,14937 ,16434 ,24189 ,4786 ,20299 ,1494 ,15463 ,2801 ,6976 ,29891 ,19337 ,27032 ,26260 ,7130 ,30457 ,28999 ,4363 ,9750 ,32095 ,8856 ,15664 ,21211 ,23939 ,5924 ,6103 ,6360 ,14661 ,13296 ,2684 ,5899 ,395 ,26142 ,29314 ,16930 ,21493 ,7925 ,30601 ,28061 ,22074 ,4512 ,10528 ,22263 ,3184 ,11348 ,25001 ,15002 ,27985 ,27765 ,14148 ,16560 ,14047 ,16103 ,23388 ,6181 ,25713 ,28468 ,19146 ,1771 ,1346 ,26255 ,24996 ,2659 ,10981 ,11118 ,30046 ,18324 ,29856 ,21929 ,7813 ,
      15578 ,17013 ,5477 ,2104 ,22790 ,9814 ,12487 ,2664 ,17187 ,19228 ,28248 ,19715 ,568 ,28797 ,10802 ,9057 ,8444 ,6726 ,10252 ,4172 ,27327 ,32196 ,17702 ,9403 ,22238 ,20531 ,32233 ,4240 ,4793 ,18134 ,16636 ,1940 ,31280 ,8073 ,13904 ,23250 ,21964 ,24348 ,18554 ,10986 ,5320 ,9908 ,25813 ,18798 ,21750 ,29732 ,20111 ,5116 ,30748 ,28749 ,12101 ,988 ,7030 ,13999 ,31318 ,5497 ,22049 ,30609 ,27202 ,12334 ,7708 ,3729 ,16908 ,148 ,8182 ,14777 ,23163 ,2158 ,21849 ,12973 ,3082 ,11123 ,29631 ,26687 ,24817 ,10893 ,7361 ,1546 ,18921 ,20410 ,19112 ,23689 ,2212 ,2576 ,10122 ,9525 ,4138 ,2124 ,16078 ,20986 ,2459 ,11230 ,170 ,3401 ,26845 ,7700 ,28663 ,31726 ,22723 ,11643 ,30858 ,16209 ,14712 ,30051 ,6002 ,10723 ,1126 ,6205 ,24493 ,22875 ,16755 ,26429 ,30772 ,5649 ,21406 ,18262 ,31218 ,30796 ,24904 ,21089 ,14123 ,22626 ,13600 ,15658 ,9051 ,20404 ,24069 ,532 ,10447 ,5095 ,4891 ,31672 ,7848 ,12149 ,3005 ,18329 ,3504 ,2299 ,18406 ,26977 ,17618 ,6805 ,763 ,24075 ,9589 ,24751 ,30943 ,5252 ,29416 ,343 ,19490 ,17033 ,6156 ,8219 ,9178 ,8268 ,20306 ,26535 ,13472 ,16411 ,30571 ,26112 ,14631 ,21181 ,4333 ,8826 ,15433 ,29861 ,24966 ,28438 ,29826 ,2629 ,10498 ,11318 ,27955 ,16530 ,13576 ,15853 ,7475 ,10156 ,23464 ,28084 ,31413 ,3913 ,1321 ,24655 ,28686 ,24592 ,652 ,21624 ,1933 ,16404 ,118 ,27172 ,13969 ,30718 ,18768 ,20081 ,8043 ,21934 ,9373 ,10222 ,18104 ,22208 ,2074 ,12457 ,19198 ,538 ,26399 ,1096 ,16179 ,28633 ,15628 ,24039 ,5619 ,31188 ,11093 ,23133 ,1516 ,29601 ,2546 ,4108 ,20956 ,140 ,16381 ,9148 ,313 ,9559 ,26947 ,733 ,5065 ,7818 ,3883 ,7445 ,21594 ,1291 ,21151 ,15403 ,28408 ,10468 ,508 ,18074 ,20051 ,88 ,29571 ,20926 ,1066 ,15598 ,7788 ,283 ,15373 ,3853 ,58 ,1036 ,253 ,28 ,
      238 ,1021 ,7773 ,3838 ,20036 ,18059 ,29556 ,15583 ,5050 ,718 ,16366 ,9544 ,21579 ,7430 ,21136 ,10453 ,19183 ,12442 ,9358 ,22193 ,13954 ,27157 ,18753 ,21919 ,5604 ,24024 ,26384 ,28618 ,1501 ,23118 ,2531 ,125 ,13457 ,26520 ,6141 ,8253 ,30928 ,24736 ,29401 ,17018 ,2990 ,12134 ,10432 ,31657 ,18391 ,2284 ,17603 ,24060 ,27940 ,11303 ,24951 ,2614 ,14616 ,26097 ,4318 ,29846 ,31398 ,28069 ,13561 ,10141 ,28671 ,24640 ,637 ,16389 ,16893 ,3714 ,22034 ,12319 ,12086 ,28734 ,7015 ,5482 ,18539 ,24333 ,31265 ,23235 ,25798 ,9893 ,21735 ,5101 ,10787 ,28782 ,17172 ,19700 ,5462 ,16998 ,22775 ,2649 ,17687 ,32181 ,8429 ,4157 ,32218 ,20516 ,4778 ,1925 ,26830 ,3386 ,16063 ,11215 ,2197 ,23674 ,10107 ,2109 ,3067 ,12958 ,8167 ,2143 ,24802 ,26672 ,7346 ,20395 ,16740 ,22860 ,5987 ,6190 ,22708 ,31711 ,30843 ,30036 ,24889 ,30781 ,30757 ,18247 ,13585 ,22611 ,9036 ,517 ,24457 ,14188 ,6936 ,8302 ,25304 ,27537 ,5696 ,22795 ,19989 ,31351 ,13538 ,16846 ,4450 ,6448 ,4403 ,4897 ,9267 ,17876 ,19823 ,6547 ,4663 ,25169 ,2926 ,28458 ,22495 ,15788 ,12658 ,2231 ,15470 ,25585 ,10024 ,27179 ,15269 ,5530 ,9710 ,31583 ,12211 ,8962 ,29942 ,9819 ,11196 ,19681 ,3819 ,2595 ,31564 ,6528 ,14903 ,14114 ,4944 ,17523 ,6602 ,31528 ,1198 ,1369 ,29156 ,25703 ,17967 ,12848 ,30819 ,28328 ,20788 ,7918 ,26838 ,20949 ,4771 ,24174 ,21453 ,14922 ,11853 ,6245 ,25948 ,12492 ,6495 ,27504 ,10933 ,23708 ,7397 ,24703 ,20483 ,31678 ,32490 ,14333 ,13672 ,9212 ,19755 ,23741 ,20614 ,1761 ,21299 ,7063 ,27787 ,18838 ,8515 ,12036 ,24181 ,21616 ,7910 ,21478 ,5884 ,29299 ,5909 ,23924 ,6345 ,2669 ,27017 ,19322 ,1479 ,6961 ,28984 ,30442 ,9735 ,15649 ,16088 ,14032 ,14987 ,14133 ,4497 ,22059 ,22248 ,24986 ,26240 ,1331 ,6166 ,19131 ,11103 ,10966 ,18309 ,7798 ,
      23429 ,27292 ,1736 ,11716 ,23529 ,28906 ,1614 ,17192 ,25486 ,13152 ,26074 ,13820 ,32453 ,14434 ,30230 ,7854 ,8750 ,30642 ,10647 ,8981 ,25351 ,12636 ,25637 ,11338 ,27637 ,21023 ,25373 ,2478 ,2808 ,25981 ,15705 ,13976 ,869 ,18664 ,13647 ,12230 ,15116 ,20699 ,7218 ,19233 ,27584 ,11922 ,7992 ,11249 ,25885 ,21672 ,32369 ,21397 ,30124 ,15982 ,22399 ,20340 ,14550 ,12525 ,22989 ,3174 ,28522 ,22082 ,3043 ,29505 ,31734 ,31969 ,19001 ,9156 ,6066 ,12367 ,12011 ,29961 ,9660 ,11961 ,19914 ,28253 ,15964 ,11904 ,27274 ,21005 ,12922 ,11886 ,8675 ,12155 ,22842 ,12940 ,3696 ,32163 ,12424 ,700 ,26502 ,28051 ,17505 ,19663 ,14170 ,15770 ,14315 ,27486 ,21460 ,1313 ,17959 ,8693 ,21274 ,26569 ,14515 ,6278 ,22673 ,19720 ,19361 ,27235 ,3452 ,13403 ,5743 ,7529 ,19579 ,5640 ,22333 ,22342 ,30133 ,9838 ,23607 ,22966 ,12997 ,10518 ,4953 ,12173 ,26648 ,16097 ,20105 ,16749 ,27949 ,28402 ,17597 ,7340 ,14897 ,9729 ,32363 ,19573 ,32305 ,573 ,26470 ,11979 ,27917 ,3420 ,1582 ,10615 ,32337 ,3011 ,29124 ,9678 ,9992 ,13506 ,6313 ,14955 ,20451 ,27755 ,18721 ,7741 ,605 ,10400 ,6983 ,17140 ,7314 ,30725 ,8349 ,19932 ,25923 ,19027 ,8565 ,1981 ,32395 ,28802 ,13099 ,15731 ,9098 ,22139 ,30256 ,30294 ,32311 ,31209 ,23598 ,3762 ,19605 ,31602 ,5157 ,10324 ,15906 ,27975 ,8701 ,28271 ,16039 ,189 ,18429 ,21486 ,3394 ,4101 ,20509 ,12029 ,27479 ,16445 ,31032 ,24207 ,4605 ,10807 ,6884 ,16941 ,9761 ,4024 ,16571 ,13209 ,29098 ,18335 ,17785 ,10050 ,24116 ,5549 ,4429 ,25777 ,32432 ,16550 ,14235 ,29979 ,29241 ,26864 ,27349 ,16452 ,14929 ,24584 ,28320 ,181 ,7372 ,15288 ,24504 ,31101 ,1443 ,9062 ,21761 ,12385 ,24002 ,7719 ,6638 ,4804 ,579 ,21080 ,10509 ,6084 ,24275 ,663 ,23300 ,20317 ,17629 ,23378 ,11624 ,2557 ,2085 ,969 ,21162 ,5233 ,30699 ,69 ,
      11059 ,3470 ,14089 ,5286 ,5840 ,7096 ,30398 ,8449 ,4727 ,18587 ,31634 ,12771 ,24137 ,3226 ,14289 ,3510 ,25260 ,3303 ,16802 ,1388 ,12614 ,25147 ,25125 ,8846 ,17923 ,13421 ,25659 ,24836 ,29898 ,3961 ,19637 ,18775 ,21535 ,11019 ,3794 ,1217 ,9314 ,1859 ,23074 ,6731 ,27896 ,27253 ,16345 ,10912 ,17559 ,21332 ,26476 ,14703 ,22664 ,19379 ,18203 ,23323 ,8123 ,11432 ,23630 ,32085 ,18495 ,4520 ,5438 ,20225 ,22731 ,27691 ,32137 ,321 ,2764 ,3263 ,8937 ,29175 ,1692 ,13335 ,14390 ,10257 ,825 ,7547 ,21353 ,26706 ,18957 ,32644 ,15938 ,2305 ,14471 ,5761 ,13359 ,30977 ,26604 ,18871 ,22922 ,7120 ,17461 ,21997 ,28007 ,22549 ,19870 ,31039 ,11860 ,7467 ,6594 ,19597 ,15244 ,11510 ,24231 ,31461 ,5189 ,4177 ,17741 ,30191 ,24540 ,28930 ,29054 ,3593 ,11985 ,16200 ,6269 ,24381 ,10356 ,25722 ,27873 ,27561 ,19529 ,4353 ,13055 ,5658 ,28758 ,29650 ,15862 ,27820 ,28227 ,18083 ,11607 ,23283 ,28303 ,6621 ,6867 ,31015 ,17768 ,27332 ,18704 ,6296 ,17580 ,1565 ,13082 ,8548 ,23581 ,18412 ,28505 ,14533 ,852 ,25868 ,25469 ,23512 ,8733 ,2791 ,17488 ,12407 ,6049 ,12905 ,19344 ,14498 ,22316 ,20088 ,24872 ,22691 ,26813 ,24785 ,18522 ,12069 ,10770 ,32201 ,5587 ,13937 ,221 ,21562 ,2973 ,30911 ,27923 ,28654 ,17950 ,1181 ,15252 ,31547 ,19972 ,25287 ,9250 ,15453 ,21282 ,19738 ,4754 ,7380 ,27000 ,5892 ,16071 ,11086 ,17680 ,21292 ,17498 ,14228 ,17454 ,17437 ,18461 ,17707 ,17471 ,25452 ,11590 ,13065 ,5570 ,18505 ,17933 ,26983 ,18478 ,8106 ,21518 ,17542 ,4710 ,5823 ,25243 ,29881 ,17444 ,26587 ,2747 ,18940 ,17724 ,24214 ,6252 ,15845 ,17515 ,3754 ,1173 ,4963 ,18159 ,28532 ,27647 ,9408 ,25216 ,8711 ,18731 ,20429 ,14245 ,28132 ,3426 ,11634 ,26560 ,17977 ,22505 ,9623 ,21309 ,21649 ,13291 ,26250 ,17697 ,31313 ,4133 ,24899 ,19485 ,31408 ,5614 ,1061 ,
      18748 ,4313 ,22770 ,30838 ,2921 ,29151 ,20609 ,22243 ,25632 ,22984 ,26497 ,12992 ,20446 ,15901 ,32427 ,17624 ,25120 ,23625 ,22917 ,19524 ,8728 ,9245 ,25238 ,13286 ,25233 ,21783 ,28834 ,8376 ,27039 ,16251 ,13126 ,8050 ,12744 ,13015 ,6911 ,13770 ,28149 ,23810 ,8597 ,20536 ,14262 ,31930 ,31137 ,12794 ,7276 ,17812 ,1588 ,1117 ,3443 ,29765 ,2013 ,28347 ,15517 ,13843 ,21788 ,14651 ,5813 ,10536 ,16869 ,21868 ,11651 ,13705 ,11690 ,9567 ,32058 ,30151 ,6423 ,17067 ,28549 ,14366 ,31773 ,32238 ,18176 ,20144 ,19059 ,896 ,10071 ,7182 ,27611 ,6811 ,27664 ,31878 ,14831 ,12867 ,9476 ,8777 ,28839 ,21201 ,18468 ,9856 ,25513 ,3101 ,9425 ,4612 ,25955 ,23456 ,1190 ,5149 ,19964 ,17986 ,20827 ,24390 ,19388 ,4245 ,23047 ,22360 ,29774 ,11142 ,4980 ,32523 ,10621 ,10714 ,27226 ,22351 ,15991 ,27431 ,3771 ,13624 ,8381 ,6093 ,17532 ,22457 ,28710 ,14041 ,29726 ,22869 ,11312 ,15397 ,2278 ,26666 ,6522 ,30436 ,21666 ,7523 ,30288 ,4798 ,21326 ,3587 ,30905 ,28126 ,17806 ,32517 ,15090 ,769 ,13308 ,9941 ,30326 ,7937 ,2361 ,8868 ,27044 ,26132 ,2737 ,16115 ,11360 ,23182 ,26267 ,20647 ,18638 ,21941 ,22522 ,1652 ,2901 ,20807 ,1672 ,9294 ,6847 ,18139 ,11833 ,12191 ,20016 ,2177 ,9640 ,15096 ,32343 ,24484 ,5734 ,4971 ,11518 ,29450 ,17994 ,1794 ,16256 ,385 ,26577 ,5353 ,31241 ,15296 ,12705 ,29307 ,11223 ,29594 ,4150 ,18831 ,15763 ,26857 ,22542 ,18933 ,3094 ,16641 ,15217 ,16767 ,14724 ,14796 ,24916 ,19788 ,30098 ,24081 ,3566 ,20123 ,18566 ,25431 ,31330 ,24312 ,13131 ,16920 ,17714 ,17352 ,15024 ,16648 ,17270 ,10814 ,12499 ,3905 ,25695 ,27967 ,15445 ,377 ,31425 ,23774 ,23888 ,1945 ,19502 ,25846 ,22171 ,13484 ,11783 ,775 ,3017 ,26420 ,5631 ,10705 ,14759 ,20968 ,6708 ,19210 ,8055 ,30591 ,15835 ,28420 ,5077 ,8201 ,1078 ,10204 ,9130 ,265 ,
      28375 ,8010 ,1900 ,19457 ,18888 ,14679 ,16603 ,31285 ,26621 ,15045 ,21896 ,13263 ,29262 ,11473 ,20762 ,9595 ,22939 ,20564 ,13241 ,25188 ,13798 ,16824 ,12749 ,28104 ,22306 ,11267 ,10669 ,1145 ,7137 ,6378 ,12822 ,9380 ,13376 ,25080 ,8404 ,4682 ,1814 ,16300 ,20180 ,8078 ,19552 ,11940 ,18038 ,6224 ,30994 ,13314 ,29130 ,18912 ,8666 ,27602 ,26205 ,17652 ,5778 ,2702 ,13020 ,17409 ,14488 ,22271 ,18367 ,11562 ,30866 ,26768 ,31502 ,26955 ,28024 ,4273 ,16973 ,2945 ,18014 ,16321 ,28573 ,13909 ,3669 ,21690 ,1880 ,10742 ,22566 ,5942 ,11170 ,24757 ,27459 ,25903 ,1716 ,21254 ,22014 ,6121 ,6916 ,5864 ,17478 ,26793 ,14069 ,15224 ,6403 ,6891 ,6502 ,15425 ,29934 ,32387 ,10762 ,6839 ,31056 ,23957 ,924 ,23255 ,19887 ,32266 ,4056 ,23553 ,17095 ,9947 ,9684 ,1537 ,11877 ,7173 ,3129 ,28477 ,12591 ,25328 ,13775 ,23484 ,12895 ,21415 ,12110 ,6021 ,7484 ,21229 ,9793 ,20060 ,21370 ,13730 ,23210 ,19842 ,16276 ,1835 ,15179 ,21969 ,7965 ,20717 ,9335 ,22894 ,26723 ,26160 ,4637 ,30949 ,20672 ,15134 ,32571 ,797 ,7564 ,29332 ,28154 ,32616 ,842 ,4826 ,10839 ,8909 ,30464 ,3644 ,17850 ,10229 ,29478 ,7236 ,21710 ,27845 ,32661 ,413 ,31064 ,24353 ,18974 ,27716 ,15324 ,28199 ,3986 ,30332 ,9998 ,29622 ,15955 ,18167 ,24239 ,6566 ,20835 ,7609 ,23815 ,31433 ,14523 ,19251 ,29377 ,24512 ,2322 ,5917 ,2205 ,16172 ,17165 ,13665 ,3689 ,24109 ,13352 ,21511 ,14824 ,18559 ,1709 ,16669 ,16477 ,30370 ,26885 ,30509 ,24431 ,5258 ,14407 ,31994 ,16676 ,17895 ,26006 ,27088 ,8602 ,3933 ,25459 ,12248 ,2405 ,16774 ,10274 ,16948 ,27511 ,8818 ,8954 ,1973 ,12061 ,9286 ,405 ,32698 ,26311 ,10991 ,25610 ,18682 ,5028 ,26448 ,29192 ,7943 ,13512 ,10884 ,20996 ,887 ,23851 ,22636 ,3280 ,30619 ,20541 ,11404 ,2781 ,24665 ,8229 ,5410 ,23143 ,13884 ,4871 ,293 ,
      24557 ,4205 ,30011 ,12677 ,11538 ,20201 ,17314 ,5325 ,29214 ,12543 ,23095 ,16228 ,28947 ,29017 ,28958 ,29422 ,25750 ,14568 ,20740 ,11805 ,30208 ,4381 ,14267 ,15068 ,17758 ,6660 ,29678 ,2873 ,29006 ,12566 ,19296 ,18111 ,3997 ,23007 ,5962 ,2333 ,3610 ,30475 ,26734 ,9913 ,29071 ,10285 ,26896 ,18610 ,29203 ,2367 ,6319 ,23154 ,12002 ,6414 ,22577 ,2250 ,17106 ,13175 ,31935 ,7495 ,31005 ,3192 ,31374 ,30877 ,16217 ,7148 ,29273 ,741 ,23351 ,22417 ,22586 ,11755 ,31478 ,32113 ,27381 ,25818 ,24248 ,17373 ,20253 ,23860 ,30000 ,3138 ,26214 ,349 ,5206 ,6759 ,16484 ,15807 ,1245 ,20880 ,31142 ,10176 ,11597 ,20358 ,7654 ,14731 ,4194 ,9768 ,10940 ,30563 ,15261 ,8341 ,24864 ,22514 ,29470 ,10365 ,18212 ,18803 ,1416 ,16000 ,2022 ,30070 ,11527 ,8874 ,14961 ,14768 ,12358 ,30142 ,22408 ,3538 ,19614 ,15682 ,12799 ,24284 ,6611 ,8477 ,24616 ,14996 ,5314 ,5996 ,24960 ,3877 ,2984 ,3061 ,11190 ,27011 ,27578 ,19355 ,13093 ,21755 ,27890 ,17735 ,5581 ,25210 ,14256 ,23041 ,11827 ,19496 ,19546 ,19881 ,18968 ,25604 ,29065 ,1410 ,7281 ,15873 ,17570 ,29523 ,9003 ,22742 ,4370 ,29909 ,24148 ,22215 ,10373 ,9436 ,10082 ,15489 ,4991 ,32706 ,23965 ,29737 ,7287 ,22100 ,458 ,11662 ,25739 ,27050 ,20457 ,21840 ,9651 ,28540 ,31469 ,12716 ,24398 ,26278 ,17817 ,23782 ,6286 ,17281 ,24927 ,31109 ,11794 ,23932 ,23682 ,1089 ,28775 ,14326 ,12933 ,10043 ,5754 ,8099 ,31871 ,20116 ,25896 ,31987 ,6752 ,31745 ,29667 ,2819 ,32464 ,17039 ,30267 ,31752 ,30377 ,18440 ,5675 ,6994 ,1593 ,4584 ,13072 ,27360 ,16582 ,14803 ,6649 ,4031 ,23715 ,21173 ,31575 ,19019 ,24777 ,20799 ,27837 ,15481 ,4461 ,5121 ,15879 ,8526 ,7408 ,10593 ,28995 ,26138 ,27761 ,11114 ,28244 ,32229 ,25809 ,27198 ,24813 ,2455 ,1122 ,13596 ,18402 ,9174 ,29822 ,28682 ,18100 ,1512 ,21590 ,15369 ,
      16362 ,26380 ,10428 ,13557 ,31261 ,8425 ,8163 ,30753 ,13534 ,12654 ,3815 ,30815 ,10929 ,27783 ,1475 ,6162 ,26070 ,25369 ,7988 ,3039 ,27270 ,14166 ,3448 ,26644 ,27913 ,601 ,9094 ,16035 ,9757 ,29237 ,23998 ,2081 ,31630 ,25655 ,16341 ,5434 ,21349 ,28003 ,24536 ,28754 ,17576 ,6045 ,217 ,4750 ,11586 ,2743 ,18727 ,4129 ,26493 ,28830 ,31133 ,16865 ,19055 ,25509 ,29770 ,28706 ,30901 ,11356 ,20012 ,31237 ,14720 ,15020 ,22167 ,5073 ,21892 ,10665 ,18034 ,18363 ,1876 ,14065 ,4052 ,12106 ,9331 ,10835 ,15320 ,29373 ,16473 ,2401 ,5024 ,8225 ,23091 ,29674 ,26892 ,31370 ,20249 ,7650 ,2018 ,24612 ,5577 ,8999 ,454 ,24923 ,6748 ,16578 ,7404 ,29818 ,3811 ,9090 ,213 ,20008 ,15316 ,450 ,32739 ,993 ,29529 ,30660 ,32743 ,21108 ,1234 ,16121 ,7747 ,9516 ,691 ,8768 ,20871 ,19155 ,11036 ,23406 ,28352 ,27129 ,21552 ,18271 ,997 ,26356 ,10165 ,19432 ,15557 ,97 ,20368 ,25391 ,28593 ,8487 ,11449 ,3202 ,6670 ,7035 ,8140 ,17291 ,29533 ,20586 ,27370 ,31817 ,14590 ,9184 ,23647 ,19261 ,4836 ,6467 ,12258 ,3325 ,15522 ,24675 ,26803 ,2496 ,30664 ,21425 ,32102 ,22281 ,11277 ,12464 ,18220 ,17230 ,2506 ,4469 ,5373 ,26319 ,932 ,14004 ,9009 ,21041 ,32747 ,18281 ,23340 ,11366 ,611 ,19103 ,22833 ,27655 ,5197 ,7882 ,19396 ,25019 ,13848 ,23896 ,22681 ,17220 ,21112 ,1451 ,11744 ,6353 ,10115 ,15621 ,5455 ,19748 ,12417 ,4422 ,26597 ,4703 ,9469 ,31323 ,22007 ,25999 ,1238 ,5668 ,20242 ,4530 ,13431 ,8274 ,9866 ,2826 ,30516 ,22467 ,4537 ,10546 ,21793 ,25557 ,18512 ,5363 ,16125 ,19795 ,17362 ,13216 ,24710 ,28430 ,19673 ,15723 ,13929 ,12183 ,27708 ,22092 ,21033 ,5502 ,22748 ,28281 ,7751 ,14875 ,29989 ,23188 ,10406 ,2567 ,32154 ,12858 ,15798 ,4916 ,7073 ,28883 ,14656 ,1341 ,32191 ,13994 ,9520 ,30791 ,338 ,28079 ,24034 ,20921 ,
      27152 ,26092 ,16993 ,31706 ,25164 ,1364 ,23736 ,22054 ,12631 ,12520 ,695 ,22961 ,14950 ,10319 ,25772 ,20312 ,25142 ,11427 ,18866 ,27556 ,23507 ,25282 ,5818 ,21644 ,9240 ,13838 ,8772 ,13619 ,8863 ,1789 ,24307 ,19205 ,16819 ,2697 ,6116 ,25323 ,29327 ,7604 ,27083 ,30614 ,4376 ,13170 ,20875 ,15677 ,1405 ,26273 ,6989 ,2450 ,14161 ,25504 ,7645 ,23401 ,3320 ,25014 ,10541 ,28878 ,25277 ,25009 ,19159 ,26046 ,30059 ,25055 ,12293 ,7826 ,25676 ,3547 ,2259 ,5715 ,12725 ,25101 ,32039 ,27207 ,6575 ,14452 ,11040 ,22645 ,24853 ,28486 ,17661 ,26541 ,7891 ,32471 ,24438 ,4925 ,13438 ,19164 ,16874 ,16721 ,17940 ,22823 ,23410 ,30105 ,8330 ,29105 ,20490 ,10490 ,31556 ,30248 ,2965 ,9632 ,3978 ,25731 ,23332 ,12339 ,29915 ,27440 ,28356 ,8647 ,29459 ,20653 ,17146 ,20977 ,19654 ,9847 ,20349 ,22814 ,31611 ,26051 ,21873 ,672 ,31537 ,7872 ,27133 ,14142 ,18792 ,6199 ,2623 ,1285 ,31651 ,2137 ,2589 ,6955 ,11243 ,13397 ,22133 ,7713 ,10906 ,28924 ,21556 ,20423 ,12788 ,11136 ,2171 ,13478 ,6218 ,23547 ,28193 ,26442 ,18604 ,30064 ,11656 ,10587 ,4744 ,21102 ,18275 ,14869 ,15671 ,8641 ,3360 ,545 ,18811 ,1632 ,4293 ,5129 ,3243 ,10999 ,23263 ,3734 ,24154 ,5510 ,1001 ,3366 ,12347 ,18644 ,7320 ,161 ,14306 ,9416 ,4185 ,8321 ,4253 ,25060 ,13710 ,1953 ,19728 ,17210 ,26360 ,9070 ,3527 ,2677 ,2117 ,31181 ,2642 ,1754 ,28044 ,16543 ,7113 ,29874 ,21194 ,16913 ,5857 ,3926 ,10169 ,4577 ,24605 ,25550 ,16714 ,16417 ,30415 ,17046 ,5265 ,14207 ,8281 ,12298 ,11695 ,16424 ,26990 ,11734 ,19436 ,24088 ,8466 ,18342 ,31685 ,16522 ,14106 ,31201 ,28646 ,24476 ,29614 ,21832 ,19095 ,153 ,22221 ,27310 ,15561 ,551 ,5303 ,21947 ,30731 ,7691 ,1304 ,23447 ,30554 ,10481 ,3487 ,7831 ,9572 ,20289 ,11076 ,15611 ,101 ,2057 ,3866 ,26930 ,491 ,41 ,
      20894 ,9116 ,4076 ,10190 ,8794 ,15821 ,6773 ,8187 ,9493 ,14745 ,20372 ,10691 ,9782 ,6694 ,29700 ,30577 ,28856 ,23874 ,17387 ,23760 ,3152 ,25681 ,32063 ,363 ,32127 ,22157 ,25395 ,25832 ,21218 ,11769 ,22431 ,26406 ,14848 ,30084 ,16014 ,19774 ,8888 ,15203 ,2852 ,14782 ,10379 ,15749 ,28597 ,18817 ,12884 ,22528 ,8355 ,16627 ,15696 ,13117 ,19287 ,24298 ,31895 ,3552 ,30156 ,25417 ,27681 ,15010 ,8491 ,17338 ,6010 ,17256 ,27405 ,3891 ,25530 ,18624 ,10299 ,20633 ,2381 ,2723 ,31797 ,23168 ,30489 ,30312 ,11453 ,9927 ,3118 ,2347 ,23021 ,26118 ,13189 ,30274 ,14414 ,7509 ,9873 ,2264 ,6428 ,30422 ,18485 ,30891 ,3206 ,3573 ,7162 ,17792 ,32497 ,755 ,4395 ,32329 ,23573 ,15082 ,4629 ,11819 ,14582 ,2163 ,9442 ,2887 ,6674 ,1638 ,12580 ,1658 ,19938 ,18125 ,25972 ,16242 ,12557 ,1780 ,29031 ,5720 ,17072 ,29436 ,20215 ,31227 ,7039 ,5339 ,23473 ,12691 ,4219 ,29580 ,19076 ,11676 ,22114 ,13691 ,27064 ,5799 ,32020 ,21854 ,32720 ,1999 ,8144 ,29751 ,913 ,15503 ,9450 ,14637 ,26292 ,8583 ,15160 ,23796 ,20161 ,12730 ,28554 ,13756 ,18193 ,31123 ,17295 ,31916 ,23946 ,7262 ,31852 ,1103 ,1424 ,32413 ,32286 ,15887 ,7199 ,25618 ,19895 ,12978 ,10088 ,22756 ,29537 ,4299 ,29923 ,2907 ,25929 ,22229 ,27628 ,25224 ,17749 ,9231 ,23055 ,25106 ,14371 ,19510 ,19369 ,28820 ,20590 ,21769 ,6828 ,27025 ,3075 ,8036 ,7008 ,25941 ,19907 ,4598 ,14383 ,18454 ,31766 ,3087 ,28566 ,14817 ,27374 ,31864 ,4045 ,9462 ,32032 ,21187 ,31790 ,31759 ,32001 ,14352 ,2833 ,32044 ,31778 ,17053 ,8113 ,19045 ,31821 ,20130 ,32255 ,10057 ,14340 ,6797 ,6440 ,10607 ,8540 ,32509 ,26152 ,23033 ,31809 ,11128 ,15495 ,19950 ,14594 ,5135 ,17084 ,20813 ,19033 ,4231 ,2469 ,8367 ,2864 ,13610 ,30168 ,27212 ,32243 ,27417 ,32075 ,28696 ,9188 ,22443 ,1526 ,29712 ,6785 ,15383 ,
      29791 ,28213 ,27730 ,27806 ,30346 ,13041 ,31840 ,29636 ,427 ,10342 ,23651 ,24367 ,11159 ,27859 ,7250 ,4339 ,7623 ,5175 ,26183 ,31447 ,22377 ,6580 ,18181 ,11496 ,23064 ,24526 ,19265 ,30177 ,5931 ,29040 ,31904 ,16186 ,29346 ,15924 ,9967 ,32630 ,32540 ,811 ,15148 ,26692 ,4997 ,8923 ,4840 ,3249 ,3658 ,1678 ,8571 ,10243 ,10638 ,22908 ,20731 ,18857 ,26174 ,14457 ,20149 ,30963 ,1849 ,27993 ,6471 ,21983 ,10731 ,19856 ,13744 ,7453 ,27102 ,19623 ,17115 ,3947 ,24407 ,17909 ,32008 ,24822 ,20844 ,16788 ,12262 ,3289 ,16962 ,12600 ,5787 ,8832 ,19405 ,30384 ,16683 ,7082 ,30523 ,11045 ,19064 ,5272 ,21525 ,31620 ,3329 ,18573 ,4262 ,24123 ,13679 ,3496 ,19981 ,26462 ,18696 ,21318 ,7957 ,27882 ,8132 ,10898 ,32712 ,3780 ,15526 ,11005 ,18003 ,9300 ,1987 ,6717 ,30633 ,23616 ,14559 ,11418 ,5166 ,22650 ,901 ,23309 ,1207 ,5424 ,24679 ,4506 ,13898 ,22717 ,14625 ,307 ,6135 ,16057 ,9704 ,5878 ,13641 ,21268 ,25917 ,7366 ,3788 ,15238 ,26807 ,1167 ,6905 ,19958 ,2895 ,15439 ,8398 ,10756 ,21704 ,12055 ,5956 ,24858 ,10076 ,24771 ,16335 ,207 ,2500 ,13923 ,6110 ,2959 ,4287 ,28640 ,16008 ,23567 ,32280 ,8534 ,9961 ,18690 ,32274 ,1551 ,23971 ,28289 ,30668 ,23269 ,27448 ,6853 ,32401 ,27318 ,25342 ,8719 ,30199 ,23498 ,22368 ,28491 ,7187 ,25854 ,27243 ,6035 ,21429 ,12393 ,21243 ,19330 ,12966 ,20074 ,28727 ,6238 ,11954 ,24200 ,13328 ,17430 ,14359 ,18926 ,16314 ,21504 ,32106 ,8092 ,14058 ,4696 ,25094 ,29867 ,2716 ,18447 ,17902 ,17423 ,22474 ,17666 ,27616 ,14214 ,17549 ,11576 ,22285 ,25438 ,26782 ,5556 ,9219 ,26969 ,16838 ,3412 ,1557 ,28118 ,22886 ,25202 ,20578 ,20415 ,29743 ,1159 ,11281 ,3740 ,6392 ,18145 ,28808 ,9394 ,11329 ,13277 ,15059 ,21635 ,11487 ,26546 ,6816 ,9609 ,14693 ,4119 ,12468 ,31299 ,15414 ,19471 ,8024 ,1047 ,
      31154 ,18295 ,21055 ,10952 ,11380 ,26226 ,27393 ,19117 ,26333 ,14973 ,18224 ,14018 ,12811 ,4483 ,17244 ,24972 ,25033 ,6331 ,26746 ,23910 ,31947 ,7896 ,27669 ,29285 ,14279 ,1465 ,17234 ,19308 ,6367 ,28970 ,17326 ,15635 ,3339 ,20469 ,23977 ,24689 ,17829 ,6481 ,19275 ,23694 ,7293 ,21439 ,2510 ,24160 ,22295 ,11839 ,13105 ,12478 ,1605 ,20600 ,17305 ,23727 ,31831 ,32476 ,31883 ,9198 ,3216 ,27773 ,4473 ,7049 ,1134 ,8501 ,25405 ,21602 ,10560 ,10010 ,31076 ,25571 ,23827 ,22481 ,2840 ,2217 ,28166 ,19809 ,5377 ,17862 ,13230 ,4649 ,15191 ,28444 ,8614 ,5682 ,26013 ,27523 ,4544 ,24443 ,14836 ,8288 ,4717 ,13524 ,26323 ,31337 ,20553 ,4436 ,19762 ,4883 ,6928 ,14889 ,28295 ,6514 ,23202 ,11182 ,28585 ,2581 ,22106 ,9696 ,936 ,5516 ,13787 ,12197 ,15737 ,9805 ,28897 ,29142 ,20192 ,1355 ,13032 ,4930 ,12872 ,31514 ,12761 ,30805 ,14008 ,12834 ,28093 ,20774 ,16615 ,20935 ,7664 ,623 ,944 ,24626 ,13860 ,31384 ,29688 ,10127 ,15534 ,24937 ,9013 ,11289 ,16592 ,14602 ,6682 ,29832 ,21805 ,29387 ,10849 ,24722 ,2415 ,13443 ,9481 ,8239 ,14079 ,10418 ,21045 ,12120 ,14668 ,18377 ,10679 ,24046 ,2030 ,21122 ,30674 ,7416 ,16135 ,5036 ,4064 ,9530 ,464 ,7759 ,32751 ,1007 ,28364 ,20022 ,9104 ,15569 ,23420 ,18739 ,24548 ,27143 ,29782 ,19169 ,8782 ,22179 ,3460 ,26370 ,18285 ,24010 ,19446 ,1487 ,8175 ,111 ,16886 ,4764 ,6059 ,20502 ,2757 ,17673 ,32051 ,4143 ,28017 ,17158 ,23344 ,28768 ,21885 ,5448 ,25669 ,2635 ,25523 ,7001 ,27095 ,28720 ,10553 ,16879 ,28844 ,12305 ,5830 ,31251 ,11370 ,24319 ,15034 ,25784 ,23748 ,5087 ,14180 ,7332 ,23275 ,26658 ,13722 ,3053 ,25383 ,2129 ,11668 ,16049 ,615 ,3372 ,29251 ,2183 ,22145 ,2095 ,11707 ,30829 ,12668 ,31697 ,27797 ,16726 ,21206 ,6176 ,8439 ,30743 ,19107 ,30767 ,9584 ,13571 ,26394 ,503 ,
      19178 ,27935 ,10782 ,16735 ,9262 ,4939 ,32485 ,16083 ,8745 ,30119 ,22837 ,22328 ,29119 ,23593 ,17780 ,10504 ,25255 ,22659 ,14466 ,6264 ,28500 ,17945 ,18473 ,26555 ,25115 ,3438 ,27659 ,27221 ,13303 ,5729 ,3561 ,5626 ,22934 ,8661 ,27454 ,11872 ,20667 ,15950 ,14402 ,20991 ,25745 ,11997 ,5201 ,12353 ,19541 ,9646 ,30262 ,28239 ,26065 ,26488 ,23086 ,686 ,23642 ,22828 ,9861 ,32149 ,25137 ,14156 ,7886 ,19649 ,6213 ,14301 ,30410 ,1299 ,28851 ,15691 ,13184 ,25967 ,26287 ,27623 ,31785 ,2464 ,7618 ,10633 ,19400 ,30628 ,8393 ,25337 ,2711 ,11324 ,25028 ,1600 ,8609 ,28892 ,21800 ,23415 ,25518 ,11702 ,25250 ,26060 ,25023 ,13138 ,25069 ,32439 ,20621 ,7840 ,25296 ,32355 ,6859 ,21658 ,16268 ,27570 ,11441 ,11235 ,27056 ,13633 ,13852 ,18650 ,1803 ,15102 ,30300 ,19219 ,13143 ,22975 ,12534 ,12511 ,10333 ,30110 ,3106 ,20326 ,1378 ,3029 ,23900 ,22068 ,8067 ,31720 ,26106 ,9142 ,26514 ,3380 ,5524 ,21472 ,18658 ,8687 ,19926 ,175 ,11013 ,19591 ,22685 ,3748 ,13009 ,5143 ,1646 ,27961 ,25074 ,32381 ,7230 ,1967 ,23001 ,8335 ,9430 ,19013 ,25649 ,9084 ,17224 ,15717 ,2691 ,30242 ,1626 ,31195 ,30078 ,32323 ,32407 ,10601 ,15918 ,26456 ,23561 ,3406 ,20463 ,14883 ,21116 ,7326 ,8655 ,32349 ,32317 ,559 ,32444 ,20437 ,28938 ,14941 ,11150 ,29110 ,4617 ,13492 ,13411 ,591 ,1455 ,7727 ,17641 ,6969 ,2151 ,30711 ,12312 ,14915 ,29954 ,16438 ,29168 ,14221 ,17060 ,26850 ,2938 ,24102 ,11748 ,10036 ,18356 ,4415 ,5708 ,16536 ,20626 ,4591 ,3940 ,24193 ,25564 ,20495 ,25960 ,16431 ,29888 ,9747 ,6357 ,16927 ,22260 ,16557 ,1768 ,18321 ,22787 ,565 ,27324 ,4790 ,21961 ,21747 ,7027 ,7705 ,21846 ,7358 ,10119 ,167 ,30855 ,24490 ,31215 ,9048 ,7845 ,17615 ,29413 ,20303 ,4330 ,10495 ,23461 ,649 ,18765 ,2071 ,15625 ,2543 ,26944 ,21148 ,29568 ,55 ,
      20033 ,21576 ,13951 ,1498 ,30925 ,18388 ,14613 ,28668 ,12083 ,25795 ,5459 ,32215 ,2194 ,24799 ,22705 ,13582 ,25301 ,4447 ,4660 ,15467 ,12208 ,31561 ,1195 ,20785 ,11850 ,7394 ,19752 ,8512 ,5906 ,28981 ,4494 ,11100 ,23526 ,32450 ,25348 ,2805 ,15113 ,25882 ,14547 ,31731 ,9657 ,12919 ,12421 ,14312 ,14512 ,5740 ,23604 ,20102 ,32360 ,1579 ,6310 ,6980 ,8562 ,30253 ,5154 ,18426 ,31029 ,16568 ,4426 ,27346 ,24501 ,6635 ,23297 ,21159 ,5837 ,24134 ,12611 ,29895 ,9311 ,17556 ,8120 ,22728 ,1689 ,18954 ,26601 ,19867 ,24228 ,29051 ,27870 ,15859 ,6864 ,13079 ,25466 ,19341 ,18519 ,2970 ,19969 ,26997 ,17451 ,5567 ,4707 ,17721 ,18156 ,14242 ,21306 ,19482 ,2918 ,20443 ,8725 ,27036 ,28146 ,7273 ,15514 ,11648 ,28546 ,10068 ,9473 ,9422 ,20824 ,4977 ,3768 ,29723 ,21663 ,17803 ,2358 ,26264 ,1669 ,9637 ,17991 ,12702 ,22539 ,24913 ,31327 ,17267 ,31422 ,11780 ,6705 ,1075 ,18885 ,29259 ,13795 ,7134 ,1811 ,30991 ,5775 ,30863 ,18011 ,22563 ,22011 ,6400 ,31053 ,17092 ,12588 ,7481 ,16273 ,26720 ,7561 ,30461 ,32658 ,3983 ,20832 ,2319 ,13349 ,26882 ,26003 ,10271 ,402 ,29189 ,3277 ,23140 ,11535 ,28944 ,30205 ,29003 ,3607 ,29200 ,17103 ,16214 ,31475 ,29997 ,1242 ,4191 ,29467 ,11524 ,19611 ,5311 ,27575 ,14253 ,29062 ,4367 ,4988 ,25736 ,24395 ,11791 ,5751 ,29664 ,5672 ,6646 ,27834 ,28992 ,24810 ,18097 ,31258 ,10926 ,27267 ,9754 ,21346 ,11583 ,19052 ,14717 ,1873 ,16470 ,20246 ,6745 ,15313 ,1231 ,11033 ,10162 ,11446 ,27367 ,12255 ,32099 ,5370 ,23337 ,19393 ,11741 ,26594 ,20239 ,4534 ,17359 ,27705 ,29986 ,7070 ,335 ,25161 ,14947 ,23504 ,8860 ,29324 ,1402 ,3317 ,30056 ,12722 ,24850 ,13435 ,8327 ,3975 ,29456 ,31608 ,18789 ,11240 ,12785 ,18601 ,15668 ,3240 ,12344 ,4250 ,3524 ,7110 ,24602 ,8278 ,8463 ,29611 ,5300 ,3484 ,3863 ,
      8791 ,9779 ,3149 ,21215 ,8885 ,12881 ,31892 ,6007 ,2378 ,3115 ,9870 ,7159 ,4626 ,12577 ,29028 ,23470 ,27061 ,910 ,20158 ,23943 ,7196 ,29920 ,23052 ,6825 ,14380 ,4042 ,2830 ,32252 ,26149 ,17081 ,30165 ,1523 ,30343 ,11156 ,22374 ,5928 ,32537 ,3655 ,26171 ,10728 ,24404 ,16959 ,30520 ,4259 ,7954 ,18000 ,5163 ,13895 ,13638 ,6902 ,5953 ,6107 ,9958 ,27445 ,22365 ,21240 ,13325 ,14055 ,22471 ,26779 ,22883 ,6389 ,11484 ,15411 ,11377 ,12808 ,31944 ,6364 ,17826 ,22292 ,31828 ,1131 ,23824 ,13227 ,4541 ,20550 ,23199 ,13784 ,13029 ,28090 ,13857 ,16589 ,2412 ,14665 ,16132 ,28361 ,29779 ,19443 ,2754 ,21882 ,10550 ,15031 ,13719 ,29248 ,27794 ,9581 ,9259 ,29116 ,28497 ,13300 ,20664 ,19538 ,23639 ,6210 ,26284 ,8390 ,21797 ,25066 ,16265 ,1800 ,10330 ,8064 ,18655 ,13006 ,22998 ,2688 ,15915 ,8652 ,11147 ,17638 ,29165 ,18353 ,25561 ,22257 ,21958 ,30852 ,4327 ,26941 ,30922 ,2191 ,12205 ,5903 ,15110 ,14509 ,8559 ,24498 ,9308 ,24225 ,18516 ,18153 ,28143 ,20821 ,1666 ,31419 ,1808 ,31050 ,32655 ,399 ,3604 ,29464 ,4985 ,27831 ,21343 ,15310 ,5367 ,27702 ,29321 ,3972 ,3237 ,29608 ,8882 ,4623 ,7193 ,26146 ,32534 ,7951 ,9955 ,22880 ,17823 ,23196 ,16129 ,13716 ,20661 ,16262 ,15912 ,21955 ,15107 ,28140 ,3601 ,29318 ,32531 ,20658 ,32528 ,783 ,7537 ,10825 ,19799 ,4812 ,786 ,30450 ,26680 ,10215 ,24326 ,27497 ,11897 ,16934 ,7540 ,25445 ,20137 ,16760 ,21683 ,16662 ,17366 ,31980 ,10828 ,25992 ,14445 ,3919 ,30305 ,14810 ,16781 ,21497 ,19802 ,17151 ,10626 ,24095 ,18947 ,16463 ,13220 ,16655 ,4815 ,26871 ,18845 ,5244 ,6539 ,13498 ,25860 ,7929 ,789 ,25596 ,6459 ,26434 ,23788 ,12047 ,24714 ,1959 ,30453 ,391 ,27981 ,10977 ,19224 ,20527 ,9904 ,30605 ,26683 ,20982 ,10719 ,22622 ,2295 ,8215 ,28434 ,24651 ,10218 ,23129 ,7441 ,279 ,
      714 ,24020 ,12130 ,28065 ,24329 ,32177 ,12954 ,30777 ,31347 ,15784 ,19677 ,12844 ,27500 ,7059 ,19318 ,1327 ,13148 ,21019 ,11918 ,22078 ,11900 ,19659 ,27231 ,12169 ,11975 ,7737 ,15727 ,28267 ,16937 ,29975 ,12381 ,2553 ,18583 ,13417 ,27249 ,4516 ,7543 ,21993 ,30187 ,5654 ,6292 ,12403 ,13933 ,19734 ,25448 ,26583 ,8707 ,31309 ,22980 ,21779 ,31926 ,10532 ,20140 ,9852 ,22356 ,22453 ,3583 ,16111 ,12187 ,5349 ,16763 ,17348 ,25842 ,28416 ,15041 ,11263 ,11936 ,22267 ,21686 ,26789 ,32262 ,21411 ,20713 ,4822 ,27712 ,19247 ,16665 ,12244 ,18678 ,24661 ,12539 ,6656 ,10281 ,3188 ,17369 ,20354 ,15996 ,8473 ,17731 ,29519 ,22096 ,17277 ,31983 ,27356 ,8522 ,9170 ,12650 ,597 ,6041 ,11352 ,10831 ,8995 ,30656 ,18267 ,17287 ,2492 ,21037 ,17216 ,25995 ,5359 ,28277 ,13990 ,12516 ,13834 ,13166 ,25005 ,14448 ,22819 ,27436 ,7868 ,28920 ,21098 ,5506 ,17206 ,3922 ,11730 ,27306 ,15607 ,14741 ,22153 ,15745 ,15006 ,30308 ,30887 ,2883 ,31223 ,1995 ,31119 ,22752 ,28816 ,14813 ,19041 ,19946 ,28692 ,10338 ,24522 ,8919 ,27989 ,16784 ,31616 ,3776 ,5420 ,15234 ,203 ,28285 ,6031 ,21500 ,11572 ,1155 ,4115 ,14969 ,1461 ,21435 ,27769 ,19805 ,13520 ,9692 ,30801 ,24933 ,10414 ,7755 ,26366 ,17154 ,31247 ,16045 ,30739 ,30115 ,3434 ,11993 ,14152 ,10629 ,26056 ,13629 ,3025 ,19587 ,9080 ,14879 ,587 ,24098 ,9743 ,7354 ,2067 ,25791 ,7390 ,12915 ,16564 ,18950 ,5563 ,10064 ,24909 ,22559 ,26878 ,29993 ,29660 ,16466 ,20235 ,24846 ,24598 ,3111 ,4038 ,16955 ,14051 ,13223 ,21878 ,8386 ,18349 ,24221 ,15306 ,23192 ,10821 ,16658 ,16459 ,12043 ,8211 ,15780 ,7733 ,12399 ,16107 ,4818 ,29515 ,2488 ,21094 ,31115 ,199 ,10410 ,9076 ,26874 ,15302 ,195 ,979 ,20331 ,28338 ,2241 ,23392 ,18848 ,677 ,6098 ,19141 ,4167 ,983 ,2571 ,18257 ,5247 ,10151 ,28628 ,83 ,
      22188 ,2609 ,19695 ,6185 ,6542 ,31523 ,9207 ,14128 ,8976 ,20335 ,32158 ,9833 ,13501 ,31597 ,5544 ,658 ,1383 ,23318 ,30972 ,25717 ,25863 ,31542 ,17537 ,9618 ,19519 ,28342 ,12862 ,27426 ,7932 ,29445 ,25426 ,20963 ,25183 ,17647 ,21249 ,28472 ,792 ,6561 ,17890 ,22631 ,11800 ,2245 ,15802 ,3533 ,25599 ,12711 ,18435 ,27193 ,3034 ,16860 ,31365 ,19150 ,6462 ,7877 ,22462 ,4911 ,27551 ,23396 ,4920 ,22809 ,26437 ,8316 ,14202 ,10476 ,23755 ,24293 ,7504 ,1775 ,23791 ,9226 ,14347 ,13605 ,31442 ,18852 ,7077 ,11413 ,12050 ,23493 ,17418 ,21630 ,23905 ,23722 ,27518 ,1350 ,24717 ,27138 ,28715 ,31692 ,6259 ,681 ,28887 ,12506 ,1962 ,14936 ,24188 ,20298 ,15462 ,6975 ,19336 ,26259 ,30456 ,4362 ,32094 ,15663 ,23938 ,6102 ,14660 ,2683 ,394 ,29313 ,21492 ,30600 ,22073 ,10527 ,3183 ,25000 ,27984 ,14147 ,14046 ,23387 ,25712 ,19145 ,1345 ,24995 ,10980 ,30045 ,29855 ,7812 ,17012 ,2103 ,9813 ,2663 ,19227 ,19714 ,28796 ,9056 ,6725 ,4171 ,32195 ,9402 ,20530 ,4239 ,18133 ,1939 ,8072 ,23249 ,24347 ,10985 ,9907 ,18797 ,29731 ,5115 ,28748 ,987 ,13998 ,5496 ,30608 ,12333 ,3728 ,147 ,14776 ,2157 ,12972 ,11122 ,26686 ,10892 ,1545 ,20409 ,23688 ,2575 ,9524 ,2123 ,20985 ,11229 ,3400 ,7699 ,31725 ,11642 ,16208 ,30050 ,10722 ,6204 ,22874 ,26428 ,5648 ,18261 ,30795 ,21088 ,22625 ,15657 ,20403 ,531 ,5094 ,31671 ,12148 ,18328 ,2298 ,26976 ,6804 ,24074 ,24750 ,5251 ,342 ,17032 ,8218 ,8267 ,26534 ,16410 ,26111 ,21180 ,8825 ,29860 ,28437 ,2628 ,11317 ,16529 ,15852 ,10155 ,28083 ,3912 ,24654 ,24591 ,21623 ,16403 ,27171 ,30717 ,20080 ,21933 ,10221 ,22207 ,12456 ,537 ,1095 ,28632 ,24038 ,31187 ,23132 ,29600 ,4107 ,139 ,9147 ,9558 ,732 ,7817 ,7444 ,1290 ,15402 ,10467 ,18073 ,87 ,20925 ,15597 ,282 ,3852 ,1035 ,27 ,
      1020 ,3837 ,18058 ,15582 ,717 ,9543 ,7429 ,10452 ,12441 ,22192 ,27156 ,21918 ,24023 ,28617 ,23117 ,124 ,26519 ,8252 ,24735 ,17017 ,12133 ,31656 ,2283 ,24059 ,11302 ,2613 ,26096 ,29845 ,28068 ,10140 ,24639 ,16388 ,3713 ,12318 ,28733 ,5481 ,24332 ,23234 ,9892 ,5100 ,28781 ,19699 ,16997 ,2648 ,32180 ,4156 ,20515 ,1924 ,3385 ,11214 ,23673 ,2108 ,12957 ,2142 ,26671 ,20394 ,22859 ,6189 ,31710 ,30035 ,30780 ,18246 ,22610 ,516 ,14187 ,8301 ,27536 ,22794 ,31350 ,16845 ,6447 ,4896 ,17875 ,6546 ,25168 ,28457 ,15787 ,2230 ,25584 ,27178 ,5529 ,31582 ,8961 ,9818 ,19680 ,2594 ,6527 ,14113 ,17522 ,31527 ,1368 ,25702 ,12847 ,28327 ,7917 ,20948 ,24173 ,14921 ,6244 ,12491 ,27503 ,23707 ,24702 ,31677 ,14332 ,9211 ,23740 ,1760 ,7062 ,18837 ,12035 ,21615 ,21477 ,29298 ,23923 ,2668 ,19321 ,6960 ,30441 ,15648 ,14031 ,14132 ,22058 ,24985 ,1330 ,19130 ,10965 ,7797 ,27291 ,11715 ,28905 ,17191 ,13151 ,13819 ,14433 ,7853 ,30641 ,8980 ,12635 ,11337 ,21022 ,2477 ,25980 ,13975 ,18663 ,12229 ,20698 ,19232 ,11921 ,11248 ,21671 ,21396 ,15981 ,20339 ,12524 ,3173 ,22081 ,29504 ,31968 ,9155 ,12366 ,29960 ,11960 ,28252 ,11903 ,21004 ,11885 ,12154 ,12939 ,32162 ,699 ,28050 ,19662 ,15769 ,27485 ,1312 ,8692 ,26568 ,6277 ,19719 ,27234 ,13402 ,7528 ,5639 ,22341 ,9837 ,22965 ,10517 ,12172 ,16096 ,16748 ,28401 ,7339 ,9728 ,19572 ,572 ,11978 ,3419 ,10614 ,3010 ,9677 ,13505 ,14954 ,27754 ,7740 ,10399 ,17139 ,30724 ,19931 ,19026 ,1980 ,28801 ,15730 ,22138 ,30293 ,31208 ,3761 ,31601 ,10323 ,27974 ,28270 ,188 ,21485 ,4100 ,12028 ,16444 ,24206 ,10806 ,16940 ,4023 ,13208 ,18334 ,10049 ,5548 ,25776 ,16549 ,29978 ,26863 ,16451 ,24583 ,180 ,15287 ,31100 ,9061 ,12384 ,7718 ,4803 ,21079 ,6083 ,662 ,20316 ,23377 ,2556 ,968 ,5232 ,68 ,
      3469 ,5285 ,7095 ,8448 ,18586 ,12770 ,3225 ,3509 ,3302 ,1387 ,25146 ,8845 ,13420 ,24835 ,3960 ,18774 ,11018 ,1216 ,1858 ,6730 ,27252 ,10911 ,21331 ,14702 ,19378 ,23322 ,11431 ,32084 ,4519 ,20224 ,27690 ,320 ,3262 ,29174 ,13334 ,10256 ,7546 ,26705 ,32643 ,2304 ,5760 ,30976 ,18870 ,7119 ,21996 ,22548 ,31038 ,7466 ,19596 ,11509 ,31460 ,4176 ,30190 ,28929 ,3592 ,16199 ,24380 ,25721 ,27560 ,4352 ,5657 ,29649 ,27819 ,18082 ,23282 ,6620 ,31014 ,27331 ,6295 ,1564 ,8547 ,18411 ,14532 ,25867 ,23511 ,2790 ,12406 ,12904 ,14497 ,20087 ,22690 ,24784 ,12068 ,32200 ,13936 ,21561 ,30910 ,28653 ,1180 ,31546 ,25286 ,15452 ,19737 ,7379 ,5891 ,11085 ,21291 ,14227 ,17436 ,17706 ,25451 ,13064 ,18504 ,26982 ,8105 ,17541 ,5822 ,29880 ,26586 ,18939 ,24213 ,15844 ,3753 ,4962 ,28531 ,9407 ,8710 ,20428 ,28131 ,11633 ,17976 ,9622 ,21648 ,26249 ,31312 ,24898 ,31407 ,1060 ,4312 ,30837 ,29150 ,22242 ,22983 ,12991 ,15900 ,17623 ,23624 ,19523 ,9244 ,13285 ,21782 ,8375 ,16250 ,8049 ,13014 ,13769 ,23809 ,20535 ,31929 ,12793 ,17811 ,1116 ,29764 ,28346 ,13842 ,14650 ,10535 ,21867 ,13704 ,9566 ,30150 ,17066 ,14365 ,32237 ,20143 ,895 ,7181 ,6810 ,31877 ,12866 ,8776 ,21200 ,9855 ,3100 ,4611 ,23455 ,5148 ,17985 ,24389 ,4244 ,22359 ,11141 ,32522 ,10713 ,22350 ,27430 ,13623 ,6092 ,22456 ,14040 ,22868 ,15396 ,26665 ,30435 ,7522 ,4797 ,3586 ,28125 ,32516 ,768 ,9940 ,7936 ,8867 ,26131 ,16114 ,23181 ,20646 ,21940 ,1651 ,20806 ,9293 ,18138 ,12190 ,2176 ,15095 ,24483 ,4970 ,29449 ,1793 ,384 ,5352 ,15295 ,29306 ,29593 ,18830 ,26856 ,18932 ,16640 ,16766 ,14795 ,19787 ,24080 ,20122 ,25430 ,24311 ,16919 ,17351 ,16647 ,10813 ,3904 ,27966 ,376 ,23773 ,1944 ,25845 ,13483 ,774 ,26419 ,10704 ,20967 ,19209 ,30590 ,28419 ,8200 ,10203 ,264 ,
      8009 ,19456 ,14678 ,31284 ,15044 ,13262 ,11472 ,9594 ,20563 ,25187 ,16823 ,28103 ,11266 ,1144 ,6377 ,9379 ,25079 ,4681 ,16299 ,8077 ,11939 ,6223 ,13313 ,18911 ,27601 ,17651 ,2701 ,17408 ,22270 ,11561 ,26767 ,26954 ,4272 ,2944 ,16320 ,13908 ,21689 ,10741 ,5941 ,24756 ,25902 ,21253 ,6120 ,5863 ,26792 ,15223 ,6890 ,15424 ,32386 ,6838 ,23956 ,23254 ,32265 ,23552 ,9946 ,1536 ,7172 ,28476 ,25327 ,23483 ,21414 ,6020 ,21228 ,20059 ,13729 ,19841 ,1834 ,21968 ,20716 ,22893 ,26159 ,30948 ,15133 ,796 ,29331 ,32615 ,4825 ,8908 ,3643 ,10228 ,7235 ,27844 ,412 ,24352 ,27715 ,28198 ,30331 ,29621 ,18166 ,6565 ,7608 ,31432 ,19250 ,24511 ,5916 ,16171 ,13664 ,24108 ,21510 ,18558 ,16668 ,30369 ,30508 ,5257 ,31993 ,17894 ,27087 ,3932 ,12247 ,16773 ,16947 ,8817 ,1972 ,9285 ,32697 ,10990 ,18681 ,26447 ,7942 ,10883 ,886 ,22635 ,30618 ,11403 ,24664 ,5409 ,13883 ,292 ,4204 ,12676 ,20200 ,5324 ,12542 ,16227 ,29016 ,29421 ,14567 ,11804 ,4380 ,15067 ,6659 ,2872 ,12565 ,18110 ,23006 ,2332 ,30474 ,9912 ,10284 ,18609 ,2366 ,23153 ,6413 ,2249 ,13174 ,7494 ,3191 ,30876 ,7147 ,740 ,22416 ,11754 ,32112 ,25817 ,17372 ,23859 ,3137 ,348 ,6758 ,15806 ,20879 ,10175 ,20357 ,14730 ,9767 ,30562 ,8340 ,22513 ,10364 ,18802 ,15999 ,30069 ,8873 ,14767 ,30141 ,3537 ,15681 ,24283 ,8476 ,14995 ,5995 ,3876 ,3060 ,27010 ,19354 ,21754 ,17734 ,25209 ,23040 ,19495 ,19880 ,25603 ,1409 ,15872 ,29522 ,22741 ,29908 ,22214 ,9435 ,15488 ,32705 ,29736 ,22099 ,11661 ,27049 ,21839 ,28539 ,12715 ,26277 ,23781 ,17280 ,31108 ,23931 ,1088 ,14325 ,10042 ,8098 ,20115 ,31986 ,31744 ,2818 ,17038 ,31751 ,18439 ,6993 ,4583 ,27359 ,14802 ,4030 ,21172 ,19018 ,20798 ,15480 ,5120 ,8525 ,10592 ,26137 ,11113 ,32228 ,27197 ,2454 ,13595 ,9173 ,28681 ,1511 ,15368 ,
      26379 ,13556 ,8424 ,30752 ,12653 ,30814 ,27782 ,6161 ,25368 ,3038 ,14165 ,26643 ,600 ,16034 ,29236 ,2080 ,25654 ,5433 ,28002 ,28753 ,6044 ,4749 ,2742 ,4128 ,28829 ,16864 ,25508 ,28705 ,11355 ,31236 ,15019 ,5072 ,10664 ,18362 ,14064 ,12105 ,10834 ,29372 ,2400 ,8224 ,29673 ,31369 ,7649 ,24611 ,8998 ,24922 ,16577 ,29817 ,9089 ,20007 ,449 ,992 ,30659 ,21107 ,16120 ,9515 ,8767 ,19154 ,23405 ,27128 ,18270 ,26355 ,19431 ,96 ,25390 ,8486 ,3201 ,7034 ,17290 ,20585 ,31816 ,9183 ,19260 ,6466 ,3324 ,24674 ,2495 ,21424 ,22280 ,12463 ,17229 ,4468 ,26318 ,14003 ,21040 ,18280 ,11365 ,19102 ,27654 ,7881 ,25018 ,23895 ,17219 ,1450 ,6352 ,15620 ,19747 ,4421 ,4702 ,31322 ,25998 ,5667 ,4529 ,8273 ,2825 ,22466 ,10545 ,25556 ,5362 ,19794 ,13215 ,28429 ,15722 ,12182 ,22091 ,5501 ,28280 ,14874 ,23187 ,2566 ,12857 ,4915 ,28882 ,1340 ,13993 ,30790 ,28078 ,20920 ,26091 ,31705 ,1363 ,22053 ,12519 ,22960 ,10318 ,20311 ,11426 ,27555 ,25281 ,21643 ,13837 ,13618 ,1788 ,19204 ,2696 ,25322 ,7603 ,30613 ,13169 ,15676 ,26272 ,2449 ,25503 ,23400 ,25013 ,28877 ,25008 ,26045 ,25054 ,7825 ,3546 ,5714 ,25100 ,27206 ,14451 ,22644 ,28485 ,26540 ,32470 ,4924 ,19163 ,16720 ,22822 ,30104 ,29104 ,10489 ,30247 ,9631 ,25730 ,12338 ,27439 ,8646 ,20652 ,20976 ,9846 ,22813 ,26050 ,671 ,7871 ,14141 ,6198 ,1284 ,2136 ,6954 ,13396 ,7712 ,28923 ,20422 ,11135 ,13477 ,23546 ,26441 ,30063 ,10586 ,21101 ,14868 ,8640 ,544 ,1631 ,5128 ,10998 ,3733 ,5509 ,3365 ,18643 ,160 ,9415 ,8320 ,25059 ,1952 ,17209 ,9069 ,2676 ,31180 ,1753 ,16542 ,29873 ,16912 ,3925 ,4576 ,25549 ,16416 ,17045 ,14206 ,12297 ,16423 ,11733 ,24087 ,18341 ,16521 ,31200 ,24475 ,21831 ,152 ,27309 ,550 ,21946 ,7690 ,23446 ,10480 ,7830 ,20288 ,15610 ,2056 ,26929 ,40 ,
      9115 ,10189 ,15820 ,8186 ,14744 ,10690 ,6693 ,30576 ,23873 ,23759 ,25680 ,362 ,22156 ,25831 ,11768 ,26405 ,30083 ,19773 ,15202 ,14781 ,15748 ,18816 ,22527 ,16626 ,13116 ,24297 ,3551 ,25416 ,15009 ,17337 ,17255 ,3890 ,18623 ,20632 ,2722 ,23167 ,30311 ,9926 ,2346 ,26117 ,30273 ,7508 ,2263 ,30421 ,30890 ,3572 ,17791 ,754 ,32328 ,15081 ,11818 ,2162 ,2886 ,1637 ,1657 ,18124 ,16241 ,1779 ,5719 ,29435 ,31226 ,5338 ,12690 ,29579 ,11675 ,13690 ,5798 ,21853 ,1998 ,29750 ,15502 ,14636 ,8582 ,23795 ,12729 ,13755 ,31122 ,31915 ,7261 ,1102 ,32412 ,15886 ,25617 ,12977 ,22755 ,4298 ,2906 ,22228 ,25223 ,9230 ,25105 ,19509 ,28819 ,21768 ,27024 ,8035 ,25940 ,4597 ,18453 ,3086 ,14816 ,31863 ,9461 ,21186 ,31758 ,14351 ,32043 ,17052 ,19044 ,20129 ,10056 ,6796 ,10606 ,32508 ,23032 ,11127 ,19949 ,5134 ,20812 ,4230 ,8366 ,13609 ,27211 ,27416 ,28695 ,22442 ,29711 ,15382 ,28212 ,27805 ,13040 ,29635 ,10341 ,24366 ,27858 ,4338 ,5174 ,31446 ,6579 ,11495 ,24525 ,30176 ,29039 ,16185 ,15923 ,32629 ,810 ,26691 ,8922 ,3248 ,1677 ,10242 ,22907 ,18856 ,14456 ,30962 ,27992 ,21982 ,19855 ,7452 ,19622 ,3946 ,17908 ,24821 ,16787 ,3288 ,12599 ,8831 ,30383 ,7081 ,11044 ,5271 ,31619 ,18572 ,24122 ,3495 ,26461 ,21317 ,27881 ,10897 ,3779 ,11004 ,9299 ,6716 ,23615 ,11417 ,22649 ,23308 ,5423 ,4505 ,22716 ,306 ,16056 ,5877 ,21267 ,7365 ,15237 ,1166 ,19957 ,15438 ,10755 ,12054 ,24857 ,24770 ,206 ,13922 ,2958 ,28639 ,23566 ,8533 ,18689 ,1550 ,28288 ,23268 ,6852 ,27317 ,8718 ,23497 ,28490 ,25853 ,6034 ,12392 ,19329 ,20073 ,6237 ,24199 ,17429 ,18925 ,21503 ,8091 ,4695 ,29866 ,18446 ,17422 ,17665 ,14213 ,11575 ,25437 ,5555 ,26968 ,3411 ,28117 ,25201 ,20414 ,1158 ,3739 ,18144 ,9393 ,13276 ,21634 ,26545 ,9608 ,4118 ,31298 ,19470 ,1046 ,
      18294 ,10951 ,26225 ,19116 ,14972 ,14017 ,4482 ,24971 ,6330 ,23909 ,7895 ,29284 ,1464 ,19307 ,28969 ,15634 ,20468 ,24688 ,6480 ,23693 ,21438 ,24159 ,11838 ,12477 ,20599 ,23726 ,32475 ,9197 ,27772 ,7048 ,8500 ,21601 ,10009 ,25570 ,22480 ,2216 ,19808 ,17861 ,4648 ,28443 ,5681 ,27522 ,24442 ,8287 ,13523 ,31336 ,4435 ,4882 ,14888 ,6513 ,11181 ,2580 ,9695 ,5515 ,12196 ,9804 ,29141 ,1354 ,4929 ,31513 ,30804 ,12833 ,20773 ,20934 ,622 ,24625 ,31383 ,10126 ,24936 ,11288 ,14601 ,29831 ,29386 ,24721 ,13442 ,8238 ,10417 ,12119 ,18376 ,24045 ,21121 ,7415 ,5035 ,9529 ,7758 ,1006 ,20021 ,15568 ,18738 ,27142 ,19168 ,22178 ,26369 ,24009 ,1486 ,110 ,4763 ,20501 ,17672 ,4142 ,17157 ,28767 ,5447 ,2634 ,7000 ,28719 ,16878 ,12304 ,31250 ,24318 ,25783 ,5086 ,7331 ,26657 ,3052 ,2128 ,16048 ,3371 ,2182 ,2094 ,30828 ,31696 ,16725 ,6175 ,30742 ,30766 ,13570 ,502 ,27934 ,16734 ,4938 ,16082 ,30118 ,22327 ,23592 ,10503 ,22658 ,6263 ,17944 ,26554 ,3437 ,27220 ,5728 ,5625 ,8660 ,11871 ,15949 ,20990 ,11996 ,12352 ,9645 ,28238 ,26487 ,685 ,22827 ,32148 ,14155 ,19648 ,14300 ,1298 ,15690 ,25966 ,27622 ,2463 ,10632 ,30627 ,25336 ,11323 ,1599 ,28891 ,23414 ,11701 ,26059 ,13137 ,32438 ,7839 ,32354 ,21657 ,27569 ,11234 ,13632 ,18649 ,15101 ,19218 ,22974 ,12510 ,30109 ,20325 ,3028 ,22067 ,31719 ,9141 ,3379 ,21471 ,8686 ,174 ,19590 ,3747 ,5142 ,27960 ,32380 ,1966 ,8334 ,19012 ,9083 ,15716 ,30241 ,31194 ,32322 ,10600 ,26455 ,3405 ,14882 ,7325 ,32348 ,558 ,20436 ,14940 ,29109 ,13491 ,590 ,7726 ,6968 ,30710 ,14914 ,16437 ,14220 ,26849 ,24101 ,10035 ,4414 ,16535 ,4590 ,24192 ,20494 ,16430 ,9746 ,16926 ,16556 ,18320 ,564 ,4789 ,21746 ,7704 ,7357 ,166 ,24489 ,9047 ,17614 ,20302 ,10494 ,648 ,2070 ,2542 ,21147 ,54 ,
      21575 ,1497 ,18387 ,28667 ,25794 ,32214 ,24798 ,13581 ,4446 ,15466 ,31560 ,20784 ,7393 ,8511 ,28980 ,11099 ,32449 ,2804 ,25881 ,31730 ,12918 ,14311 ,5739 ,20101 ,1578 ,6979 ,30252 ,18425 ,16567 ,27345 ,6634 ,21158 ,24133 ,29894 ,17555 ,22727 ,18953 ,19866 ,29050 ,15858 ,13078 ,19340 ,2969 ,26996 ,5566 ,17720 ,14241 ,19481 ,20442 ,27035 ,7272 ,11647 ,10067 ,9421 ,4976 ,29722 ,17802 ,26263 ,9636 ,12701 ,24912 ,17266 ,11779 ,1074 ,29258 ,7133 ,30990 ,30862 ,22562 ,6399 ,17091 ,7480 ,26719 ,30460 ,3982 ,2318 ,26881 ,10270 ,29188 ,23139 ,28943 ,29002 ,29199 ,16213 ,29996 ,4190 ,11523 ,5310 ,14252 ,4366 ,25735 ,11790 ,29663 ,6645 ,28991 ,18096 ,10925 ,9753 ,11582 ,14716 ,16469 ,6744 ,1230 ,10161 ,27366 ,32098 ,23336 ,11740 ,20238 ,17358 ,29985 ,334 ,14946 ,8859 ,1401 ,30055 ,24849 ,8326 ,29455 ,18788 ,12784 ,15667 ,12343 ,3523 ,24601 ,8462 ,5299 ,3862 ,9778 ,21214 ,12880 ,6006 ,3114 ,7158 ,12576 ,23469 ,909 ,23942 ,29919 ,6824 ,4041 ,32251 ,17080 ,1522 ,11155 ,5927 ,3654 ,10727 ,16958 ,4258 ,17999 ,13894 ,6901 ,6106 ,27444 ,21239 ,14054 ,26778 ,6388 ,15410 ,12807 ,6363 ,22291 ,1130 ,13226 ,20549 ,13783 ,28089 ,16588 ,14664 ,28360 ,19442 ,21881 ,15030 ,29247 ,9580 ,29115 ,13299 ,19537 ,6209 ,8389 ,25065 ,1799 ,8063 ,13005 ,2687 ,8651 ,17637 ,18352 ,22256 ,30851 ,26940 ,2190 ,5902 ,14508 ,24497 ,24224 ,18152 ,20820 ,31418 ,31049 ,398 ,29463 ,27830 ,15309 ,27701 ,3971 ,29607 ,4622 ,26145 ,7950 ,22879 ,23195 ,13715 ,16261 ,21954 ,28139 ,29317 ,20657 ,782 ,10824 ,4811 ,30449 ,10214 ,27496 ,16933 ,25444 ,16759 ,16661 ,31979 ,25991 ,3918 ,14809 ,21496 ,17150 ,24094 ,16462 ,16654 ,26870 ,5243 ,13497 ,7928 ,25595 ,26433 ,12046 ,1958 ,390 ,10976 ,20526 ,30604 ,20981 ,22621 ,8214 ,24650 ,23128 ,278 ,
      24019 ,28064 ,32176 ,30776 ,15783 ,12843 ,7058 ,1326 ,21018 ,22077 ,19658 ,12168 ,7736 ,28266 ,29974 ,2552 ,13416 ,4515 ,21992 ,5653 ,12402 ,19733 ,26582 ,31308 ,21778 ,10531 ,9851 ,22452 ,16110 ,5348 ,17347 ,28415 ,11262 ,22266 ,26788 ,21410 ,4821 ,19246 ,12243 ,24660 ,6655 ,3187 ,20353 ,8472 ,29518 ,17276 ,27355 ,9169 ,596 ,11351 ,8994 ,18266 ,2491 ,17215 ,5358 ,13989 ,13833 ,25004 ,22818 ,7867 ,21097 ,17205 ,11729 ,15606 ,22152 ,15005 ,30886 ,31222 ,31118 ,28815 ,19040 ,28691 ,24521 ,27988 ,31615 ,5419 ,202 ,6030 ,11571 ,4114 ,1460 ,27768 ,13519 ,30800 ,10413 ,26365 ,31246 ,30738 ,3433 ,14151 ,26055 ,3024 ,9079 ,586 ,9742 ,2066 ,7389 ,16563 ,5562 ,24908 ,26877 ,29659 ,20234 ,24597 ,4037 ,14050 ,21877 ,18348 ,15305 ,10820 ,16458 ,8210 ,7732 ,16106 ,29514 ,21093 ,198 ,9075 ,15301 ,978 ,28337 ,23391 ,676 ,19140 ,982 ,18256 ,10150 ,82 ,2608 ,6184 ,31522 ,14127 ,20334 ,9832 ,31596 ,657 ,23317 ,25716 ,31541 ,9617 ,28341 ,27425 ,29444 ,20962 ,17646 ,28471 ,6560 ,22630 ,2244 ,3532 ,12710 ,27192 ,16859 ,19149 ,7876 ,4910 ,23395 ,22808 ,8315 ,10475 ,24292 ,1774 ,9225 ,13604 ,18851 ,11412 ,23492 ,21629 ,23721 ,1349 ,27137 ,31691 ,680 ,12505 ,14935 ,20297 ,6974 ,26258 ,4361 ,15662 ,6101 ,2682 ,29312 ,30599 ,10526 ,24999 ,14146 ,23386 ,19144 ,24994 ,30044 ,7811 ,2102 ,2662 ,19713 ,9055 ,4170 ,9401 ,4238 ,1938 ,23248 ,10984 ,18796 ,5114 ,986 ,5495 ,12332 ,146 ,2156 ,11121 ,10891 ,20408 ,2574 ,2122 ,11228 ,7698 ,11641 ,30049 ,6203 ,26427 ,18260 ,21087 ,15656 ,530 ,31670 ,18327 ,26975 ,24073 ,5250 ,17031 ,8266 ,16409 ,21179 ,29859 ,2627 ,16528 ,10154 ,3911 ,24590 ,16402 ,30716 ,21932 ,22206 ,536 ,28631 ,31186 ,29599 ,138 ,9557 ,7816 ,1289 ,10466 ,86 ,15596 ,3851 ,26 ,
      3836 ,15581 ,9542 ,10451 ,22191 ,21917 ,28616 ,123 ,8251 ,17016 ,31655 ,24058 ,2612 ,29844 ,10139 ,16387 ,12317 ,5480 ,23233 ,5099 ,19698 ,2647 ,4155 ,1923 ,11213 ,2107 ,2141 ,20393 ,6188 ,30034 ,18245 ,515 ,8300 ,22793 ,16844 ,4895 ,6545 ,28456 ,2229 ,27177 ,31581 ,9817 ,2593 ,14112 ,31526 ,25701 ,28326 ,20947 ,14920 ,12490 ,23706 ,31676 ,9210 ,1759 ,18836 ,21614 ,29297 ,2667 ,6959 ,15647 ,14131 ,24984 ,19129 ,7796 ,11714 ,17190 ,13818 ,7852 ,8979 ,11336 ,2476 ,13974 ,12228 ,19231 ,11247 ,21395 ,20338 ,3172 ,29503 ,9154 ,29959 ,28251 ,21003 ,12153 ,32161 ,28049 ,15768 ,1311 ,26567 ,19718 ,13401 ,5638 ,9836 ,10516 ,16095 ,28400 ,9727 ,571 ,3418 ,3009 ,13504 ,27753 ,10398 ,30723 ,19025 ,28800 ,22137 ,31207 ,31600 ,27973 ,187 ,4099 ,16443 ,10805 ,4022 ,18333 ,5547 ,16548 ,26862 ,24582 ,15286 ,9060 ,7717 ,21078 ,661 ,23376 ,967 ,67 ,5284 ,8447 ,12769 ,3508 ,1386 ,8844 ,24834 ,18773 ,1215 ,6729 ,10910 ,14701 ,23321 ,32083 ,20223 ,319 ,29173 ,10255 ,26704 ,2303 ,30975 ,7118 ,22547 ,7465 ,11508 ,4175 ,28928 ,16198 ,25720 ,4351 ,29648 ,18081 ,6619 ,27330 ,1563 ,18410 ,25866 ,2789 ,12903 ,20086 ,24783 ,32199 ,21560 ,28652 ,31545 ,15451 ,7378 ,11084 ,14226 ,17705 ,13063 ,26981 ,17540 ,29879 ,18938 ,15843 ,4961 ,9406 ,20427 ,11632 ,9621 ,26248 ,24897 ,1059 ,30836 ,22241 ,12990 ,17622 ,19522 ,13284 ,8374 ,8048 ,13768 ,20534 ,12792 ,1115 ,28345 ,14649 ,21866 ,9565 ,17065 ,32236 ,894 ,6809 ,12865 ,21199 ,3099 ,23454 ,17984 ,4243 ,11140 ,10712 ,27429 ,6091 ,14039 ,15395 ,30434 ,4796 ,28124 ,767 ,7935 ,26130 ,23180 ,21939 ,20805 ,18137 ,2175 ,24482 ,29448 ,383 ,15294 ,29592 ,26855 ,16639 ,14794 ,24079 ,25429 ,16918 ,16646 ,3903 ,375 ,1943 ,13482 ,26418 ,20966 ,30589 ,8199 ,263 ,
      19455 ,31283 ,13261 ,9593 ,25186 ,28102 ,1143 ,9378 ,4680 ,8076 ,6222 ,18910 ,17650 ,17407 ,11560 ,26953 ,2943 ,13907 ,10740 ,24755 ,21252 ,5862 ,15222 ,15423 ,6837 ,23253 ,23551 ,1535 ,28475 ,23482 ,6019 ,20058 ,19840 ,21967 ,22892 ,30947 ,795 ,32614 ,8907 ,10227 ,27843 ,24351 ,28197 ,29620 ,6564 ,31431 ,24510 ,16170 ,24107 ,18557 ,30368 ,5256 ,17893 ,3931 ,16772 ,8816 ,9284 ,10989 ,26446 ,10882 ,22634 ,11402 ,5408 ,291 ,12675 ,5323 ,16226 ,29420 ,11803 ,15066 ,2871 ,18109 ,2331 ,9911 ,18608 ,23152 ,2248 ,7493 ,30875 ,739 ,11753 ,25816 ,23858 ,347 ,15805 ,10174 ,14729 ,30561 ,22512 ,18801 ,30068 ,14766 ,3536 ,24282 ,14994 ,3875 ,27009 ,21753 ,25208 ,19494 ,25602 ,15871 ,22740 ,22213 ,15487 ,29735 ,11660 ,21838 ,12714 ,23780 ,31107 ,1087 ,10041 ,20114 ,31743 ,17037 ,18438 ,4582 ,14801 ,21171 ,20797 ,5119 ,10591 ,11112 ,27196 ,13594 ,28680 ,15367 ,13555 ,30751 ,30813 ,6160 ,3037 ,26642 ,16033 ,2079 ,5432 ,28752 ,4748 ,4127 ,16863 ,28704 ,31235 ,5071 ,18361 ,12104 ,29371 ,8223 ,31368 ,24610 ,24921 ,29816 ,20006 ,991 ,21106 ,9514 ,19153 ,27127 ,26354 ,95 ,8485 ,7033 ,20584 ,9182 ,6465 ,24673 ,21423 ,12462 ,4467 ,14002 ,18279 ,19101 ,7880 ,23894 ,1449 ,15619 ,4420 ,31321 ,5666 ,8272 ,22465 ,25555 ,19793 ,28428 ,12181 ,5500 ,14873 ,2565 ,4914 ,1339 ,30789 ,20919 ,31704 ,22052 ,22959 ,20310 ,27554 ,21642 ,13617 ,19203 ,25321 ,30612 ,15675 ,2448 ,23399 ,28876 ,26044 ,7824 ,5713 ,27205 ,22643 ,26539 ,4923 ,16719 ,30103 ,10488 ,9630 ,12337 ,8645 ,20975 ,22812 ,670 ,14140 ,1283 ,6953 ,7711 ,20421 ,13476 ,26440 ,10585 ,14867 ,543 ,5127 ,3732 ,3364 ,159 ,8319 ,1951 ,9068 ,31179 ,16541 ,16911 ,4575 ,16415 ,14205 ,16422 ,24086 ,16520 ,24474 ,151 ,549 ,7689 ,10479 ,20287 ,2055 ,39 ,
      10188 ,8185 ,10689 ,30575 ,23758 ,361 ,25830 ,26404 ,19772 ,14780 ,18815 ,16625 ,24296 ,25415 ,17336 ,3889 ,20631 ,23166 ,9925 ,26116 ,7507 ,30420 ,3571 ,753 ,15080 ,2161 ,1636 ,18123 ,1778 ,29434 ,5337 ,29578 ,13689 ,21852 ,29749 ,14635 ,23794 ,13754 ,31914 ,1101 ,15885 ,12976 ,4297 ,22227 ,9229 ,19508 ,21767 ,8034 ,4596 ,3085 ,31862 ,21185 ,14350 ,17051 ,20128 ,6795 ,32507 ,11126 ,5133 ,4229 ,13608 ,27415 ,22441 ,15381 ,27804 ,29634 ,24365 ,4337 ,31445 ,11494 ,30175 ,16184 ,32628 ,26690 ,3247 ,10241 ,18855 ,30961 ,21981 ,7451 ,3945 ,24820 ,3287 ,8830 ,7080 ,5270 ,18571 ,3494 ,21316 ,10896 ,11003 ,6715 ,11416 ,23307 ,4504 ,305 ,5876 ,7364 ,1165 ,15437 ,12053 ,24769 ,13921 ,28638 ,8532 ,1549 ,23267 ,27316 ,23496 ,25852 ,12391 ,20072 ,24198 ,18924 ,8090 ,29865 ,17421 ,14212 ,25436 ,26967 ,28116 ,20413 ,3738 ,9392 ,21633 ,9607 ,31297 ,1045 ,10950 ,19115 ,14016 ,24970 ,23908 ,29283 ,19306 ,15633 ,24687 ,23692 ,24158 ,12476 ,23725 ,9196 ,7047 ,21600 ,25569 ,2215 ,17860 ,28442 ,27521 ,8286 ,31335 ,4881 ,6512 ,2579 ,5514 ,9803 ,1353 ,31512 ,12832 ,20933 ,24624 ,10125 ,11287 ,29830 ,24720 ,8237 ,12118 ,24044 ,7414 ,9528 ,1005 ,15567 ,27141 ,22177 ,24008 ,109 ,20500 ,4141 ,28766 ,2633 ,28718 ,12303 ,24317 ,5085 ,26656 ,2127 ,3370 ,2093 ,31695 ,6174 ,30765 ,501 ,16733 ,16081 ,22326 ,10502 ,6262 ,26553 ,27219 ,5624 ,11870 ,20989 ,12351 ,28237 ,684 ,32147 ,19647 ,1297 ,25965 ,2462 ,30626 ,11322 ,28890 ,11700 ,13136 ,7838 ,21656 ,11233 ,18648 ,19217 ,12509 ,20324 ,22066 ,9140 ,21470 ,173 ,3746 ,27959 ,1965 ,19011 ,15715 ,31193 ,10599 ,3404 ,7324 ,557 ,14939 ,13490 ,7725 ,30709 ,16436 ,26848 ,10034 ,16534 ,24191 ,16429 ,16925 ,18319 ,4788 ,7703 ,165 ,9046 ,20301 ,647 ,2541 ,53 ,
      1496 ,28666 ,32213 ,13580 ,15465 ,20783 ,8510 ,11098 ,2803 ,31729 ,14310 ,20100 ,6978 ,18424 ,27344 ,21157 ,29893 ,22726 ,19865 ,15857 ,19339 ,26995 ,17719 ,19480 ,27034 ,11646 ,9420 ,29721 ,26262 ,12700 ,17265 ,1073 ,7132 ,30861 ,6398 ,7479 ,30459 ,2317 ,10269 ,23138 ,29001 ,16212 ,4189 ,5309 ,4365 ,11789 ,6644 ,18095 ,9752 ,14715 ,6743 ,10160 ,32097 ,11739 ,17357 ,333 ,8858 ,30054 ,8325 ,18787 ,15666 ,3522 ,8461 ,3861 ,21213 ,6005 ,7157 ,23468 ,23941 ,6823 ,32250 ,1521 ,5926 ,10726 ,4257 ,13893 ,6105 ,21238 ,26777 ,15409 ,6362 ,1129 ,20548 ,28088 ,14663 ,19441 ,15029 ,9579 ,13298 ,6208 ,25064 ,8062 ,2686 ,17636 ,22255 ,26939 ,5901 ,24496 ,18151 ,31417 ,397 ,27829 ,27700 ,29606 ,26144 ,22878 ,13714 ,21953 ,29316 ,781 ,4810 ,10213 ,16932 ,16758 ,31978 ,3917 ,21495 ,24093 ,16653 ,5242 ,7927 ,26432 ,1957 ,10975 ,30603 ,22620 ,24649 ,277 ,28063 ,30775 ,12842 ,1325 ,22076 ,12167 ,28265 ,2551 ,4514 ,5652 ,19732 ,31307 ,10530 ,22451 ,5347 ,28414 ,22265 ,21409 ,19245 ,24659 ,3186 ,8471 ,17275 ,9168 ,11350 ,18265 ,17214 ,13988 ,25003 ,7866 ,17204 ,15605 ,15004 ,31221 ,28814 ,28690 ,27987 ,5418 ,6029 ,4113 ,27767 ,30799 ,26364 ,30737 ,14150 ,3023 ,585 ,2065 ,16562 ,24907 ,29658 ,24596 ,14049 ,18347 ,10819 ,8209 ,16105 ,21092 ,9074 ,977 ,23390 ,19139 ,18255 ,81 ,6183 ,14126 ,9831 ,656 ,25715 ,9616 ,27424 ,20961 ,28470 ,22629 ,3531 ,27191 ,19148 ,4909 ,22807 ,10474 ,1773 ,13603 ,11411 ,21628 ,1348 ,31690 ,12504 ,20296 ,26257 ,15661 ,2681 ,30598 ,24998 ,23385 ,24993 ,7810 ,2661 ,9054 ,9400 ,1937 ,10983 ,5113 ,5494 ,145 ,11120 ,20407 ,2121 ,7697 ,30048 ,26426 ,21086 ,529 ,18326 ,24072 ,17030 ,16408 ,29858 ,16527 ,3910 ,16401 ,21931 ,535 ,31185 ,137 ,7815 ,10465 ,15595 ,25 ,
      15580 ,10450 ,21916 ,122 ,17015 ,24057 ,29843 ,16386 ,5479 ,5098 ,2646 ,1922 ,2106 ,20392 ,30033 ,514 ,22792 ,4894 ,28455 ,27176 ,9816 ,14111 ,25700 ,20946 ,12489 ,31675 ,1758 ,21613 ,2666 ,15646 ,24983 ,7795 ,17189 ,7851 ,11335 ,13973 ,19230 ,21394 ,3171 ,9153 ,28250 ,12152 ,28048 ,1310 ,19717 ,5637 ,10515 ,28399 ,570 ,3008 ,27752 ,30722 ,28799 ,31206 ,27972 ,4098 ,10804 ,18332 ,16547 ,24581 ,9059 ,21077 ,23375 ,66 ,8446 ,3507 ,8843 ,18772 ,6728 ,14700 ,32082 ,318 ,10254 ,2302 ,7117 ,7464 ,4174 ,16197 ,4350 ,18080 ,27329 ,18409 ,2788 ,20085 ,32198 ,28651 ,15450 ,11083 ,17704 ,26980 ,29878 ,15842 ,9405 ,11631 ,26247 ,1058 ,22240 ,17621 ,13283 ,8047 ,20533 ,1114 ,14648 ,9564 ,32235 ,6808 ,21198 ,23453 ,4242 ,10711 ,6090 ,15394 ,4795 ,766 ,26129 ,21938 ,18136 ,24481 ,382 ,29591 ,16638 ,24078 ,16917 ,3902 ,1942 ,26417 ,30588 ,262 ,31282 ,9592 ,28101 ,9377 ,8075 ,18909 ,17406 ,26952 ,13906 ,24754 ,5861 ,15422 ,23252 ,1534 ,23481 ,20057 ,21966 ,30946 ,32613 ,10226 ,24350 ,29619 ,31430 ,16169 ,18556 ,5255 ,3930 ,8815 ,10988 ,10881 ,11401 ,290 ,5322 ,29419 ,15065 ,18108 ,9910 ,23151 ,7492 ,738 ,25815 ,346 ,10173 ,30560 ,18800 ,14765 ,24281 ,3874 ,21752 ,19493 ,15870 ,22212 ,29734 ,21837 ,23779 ,1086 ,20113 ,17036 ,4581 ,21170 ,5118 ,11111 ,13593 ,15366 ,30750 ,6159 ,26641 ,2078 ,28751 ,4126 ,28703 ,5070 ,12103 ,8222 ,24609 ,29815 ,990 ,9513 ,27126 ,94 ,7032 ,9181 ,24672 ,12461 ,14001 ,19100 ,23893 ,15618 ,31320 ,8271 ,25554 ,28427 ,5499 ,2564 ,1338 ,20918 ,22051 ,20309 ,21641 ,19202 ,30611 ,2447 ,28875 ,7823 ,27204 ,26538 ,16718 ,10487 ,12336 ,20974 ,669 ,1282 ,7710 ,13475 ,10584 ,542 ,3731 ,158 ,1950 ,31178 ,16910 ,16414 ,16421 ,16519 ,150 ,7688 ,20286 ,38 ,
      8184 ,30574 ,360 ,26403 ,14779 ,16624 ,25414 ,3888 ,23165 ,26115 ,30419 ,752 ,2160 ,18122 ,29433 ,29577 ,21851 ,14634 ,13753 ,1100 ,12975 ,22226 ,19507 ,8033 ,3084 ,21184 ,17050 ,6794 ,11125 ,4228 ,27414 ,15380 ,29633 ,4336 ,11493 ,16183 ,26689 ,10240 ,30960 ,7450 ,24819 ,8829 ,5269 ,3493 ,10895 ,6714 ,23306 ,304 ,7363 ,15436 ,24768 ,28637 ,1548 ,27315 ,25851 ,20071 ,18923 ,29864 ,14211 ,26966 ,20412 ,9391 ,9606 ,1044 ,19114 ,24969 ,29282 ,15632 ,23691 ,12475 ,9195 ,21599 ,2214 ,28441 ,8285 ,4880 ,2578 ,9802 ,31511 ,20932 ,10124 ,29829 ,8236 ,24043 ,9527 ,15566 ,22176 ,108 ,4140 ,2632 ,12302 ,5084 ,2126 ,2092 ,6173 ,500 ,16080 ,10501 ,26552 ,5623 ,20988 ,28236 ,32146 ,1296 ,2461 ,11321 ,11699 ,7837 ,11232 ,19216 ,20323 ,9139 ,172 ,27958 ,19010 ,31192 ,3403 ,556 ,13489 ,30708 ,26847 ,16533 ,16428 ,18318 ,7702 ,9045 ,646 ,52 ,28665 ,13579 ,20782 ,11097 ,31728 ,20099 ,18423 ,21156 ,22725 ,15856 ,26994 ,19479 ,11645 ,29720 ,12699 ,1072 ,30860 ,7478 ,2316 ,23137 ,16211 ,5308 ,11788 ,18094 ,14714 ,10159 ,11738 ,332 ,30053 ,18786 ,3521 ,3860 ,6004 ,23467 ,6822 ,1520 ,10725 ,13892 ,21237 ,15408 ,1128 ,28087 ,19440 ,9578 ,6207 ,8061 ,17635 ,26938 ,24495 ,31416 ,27828 ,29605 ,22877 ,21952 ,780 ,10212 ,16757 ,3916 ,24092 ,5241 ,26431 ,10974 ,22619 ,276 ,30774 ,1324 ,12166 ,2550 ,5651 ,31306 ,22450 ,28413 ,21408 ,24658 ,8470 ,9167 ,18264 ,13987 ,7865 ,15604 ,31220 ,28689 ,5417 ,4112 ,30798 ,30736 ,3022 ,2064 ,24906 ,24595 ,18346 ,8208 ,21091 ,976 ,19138 ,80 ,14125 ,655 ,9615 ,20960 ,22628 ,27190 ,4908 ,10473 ,13602 ,21627 ,31689 ,20295 ,15660 ,30597 ,23384 ,7809 ,9053 ,1936 ,5112 ,144 ,20406 ,7696 ,26425 ,528 ,24071 ,16407 ,16526 ,16400 ,534 ,136 ,10464 ,24 ,
      10449 ,121 ,24056 ,16385 ,5097 ,1921 ,20391 ,513 ,4893 ,27175 ,14110 ,20945 ,31674 ,21612 ,15645 ,7794 ,7850 ,13972 ,21393 ,9152 ,12151 ,1309 ,5636 ,28398 ,3007 ,30721 ,31205 ,4097 ,18331 ,24580 ,21076 ,65 ,3506 ,18771 ,14699 ,317 ,2301 ,7463 ,16196 ,18079 ,18408 ,20084 ,28650 ,11082 ,26979 ,15841 ,11630 ,1057 ,17620 ,8046 ,1113 ,9563 ,6807 ,23452 ,10710 ,15393 ,765 ,21937 ,24480 ,29590 ,24077 ,3901 ,26416 ,261 ,9591 ,9376 ,18908 ,26951 ,24753 ,15421 ,1533 ,20056 ,30945 ,10225 ,29618 ,16168 ,5254 ,8814 ,10880 ,289 ,29418 ,18107 ,23150 ,737 ,345 ,30559 ,14764 ,3873 ,19492 ,22211 ,21836 ,1085 ,17035 ,21169 ,11110 ,15365 ,6158 ,2077 ,4125 ,5069 ,8221 ,29814 ,9512 ,93 ,9180 ,12460 ,19099 ,15617 ,8270 ,28426 ,2563 ,20917 ,20308 ,19201 ,2446 ,7822 ,26537 ,10486 ,20973 ,1281 ,13474 ,541 ,157 ,31177 ,16413 ,16518 ,7687 ,37 ,30573 ,26402 ,16623 ,3887 ,26114 ,751 ,18121 ,29576 ,14633 ,1099 ,22225 ,8032 ,21183 ,6793 ,4227 ,15379 ,4335 ,16182 ,10239 ,7449 ,8828 ,3492 ,6713 ,303 ,15435 ,28636 ,27314 ,20070 ,29863 ,26965 ,9390 ,1043 ,24968 ,15631 ,12474 ,21598 ,28440 ,4879 ,9801 ,20931 ,29828 ,24042 ,15565 ,107 ,2631 ,5083 ,2091 ,499 ,10500 ,5622 ,28235 ,1295 ,11320 ,7836 ,19215 ,9138 ,27957 ,31191 ,555 ,30707 ,16532 ,18317 ,9044 ,51 ,13578 ,11096 ,20098 ,21155 ,15855 ,19478 ,29719 ,1071 ,7477 ,23136 ,5307 ,18093 ,10158 ,331 ,18785 ,3859 ,23466 ,1519 ,13891 ,15407 ,28086 ,9577 ,8060 ,26937 ,31415 ,29604 ,21951 ,10211 ,3915 ,5240 ,10973 ,275 ,1323 ,2549 ,31305 ,28412 ,24657 ,9166 ,13986 ,15603 ,28688 ,4111 ,30735 ,2063 ,24594 ,8207 ,975 ,79 ,654 ,20959 ,27189 ,10472 ,21626 ,20294 ,30596 ,7808 ,1935 ,143 ,7695 ,527 ,16406 ,16399 ,135 ,23 ,
      120 ,16384 ,1920 ,512 ,27174 ,20944 ,21611 ,7793 ,13971 ,9151 ,1308 ,28397 ,30720 ,4096 ,24579 ,64 ,18770 ,316 ,7462 ,18078 ,20083 ,11081 ,15840 ,1056 ,8045 ,9562 ,23451 ,15392 ,21936 ,29589 ,3900 ,260 ,9375 ,26950 ,15420 ,20055 ,10224 ,16167 ,8813 ,288 ,18106 ,736 ,30558 ,3872 ,22210 ,1084 ,21168 ,15364 ,2076 ,5068 ,29813 ,92 ,12459 ,15616 ,28425 ,20916 ,19200 ,7821 ,10485 ,1280 ,540 ,31176 ,16517 ,36 ,26401 ,3886 ,750 ,29575 ,1098 ,8031 ,6792 ,15378 ,16181 ,7448 ,3491 ,302 ,28635 ,20069 ,26964 ,1042 ,15630 ,21597 ,4878 ,20930 ,24041 ,106 ,5082 ,498 ,5621 ,1294 ,7835 ,9137 ,31190 ,30706 ,18316 ,50 ,11095 ,21154 ,19477 ,1070 ,23135 ,18092 ,330 ,3858 ,1518 ,15406 ,9576 ,26936 ,29603 ,10210 ,5239 ,274 ,2548 ,28411 ,9165 ,15602 ,4110 ,2062 ,8206 ,78 ,20958 ,10471 ,20293 ,7807 ,142 ,526 ,16398 ,22 ,16383 ,511 ,20943 ,7792 ,9150 ,28396 ,4095 ,63 ,315 ,18077 ,11080 ,1055 ,9561 ,15391 ,29588 ,259 ,26949 ,20054 ,16166 ,287 ,735 ,3871 ,1083 ,15363 ,5067 ,91 ,15615 ,20915 ,7820 ,1279 ,31175 ,35 ,3885 ,29574 ,8030 ,15377 ,7447 ,301 ,20068 ,1041 ,21596 ,20929 ,105 ,497 ,1293 ,9136 ,30705 ,49 ,21153 ,1069 ,18091 ,3857 ,15405 ,26935 ,10209 ,273 ,28410 ,15601 ,2061 ,77 ,10470 ,7806 ,525 ,21 ,510 ,7791 ,28395 ,62 ,18076 ,1054 ,15390 ,258 ,20053 ,286 ,3870 ,15362 ,90 ,20914 ,1278 ,34 ,29573 ,15376 ,300 ,1040 ,20928 ,496 ,9135 ,48 ,1068 ,3856 ,26934 ,272 ,15600 ,76 ,7805 ,20 ,7790 ,61 ,1053 ,257 ,285 ,15361 ,20913 ,33 ,15375 ,1039 ,495 ,47 ,3855 ,271 ,75 ,19 ,60 ,256 ,15360 ,32 ,1038 ,46 ,270 ,18 ,255 ,31 ,45 ,17 ,30 ,16 ,15 ,0 
   );
   constant CPIX_NORMAL_INIT_00_BIT_00_C : bit_vector(255 downto 0) := x"4F04664232E82CE1170DD0A315BB6716CFAEA193ED72F0AE40361A30FACB04F2";
   constant CPIX_NORMAL_INIT_00_BIT_01_C : bit_vector(255 downto 0) := x"467046C1196639A6E14BDE988C46CEFEDBB684FE2EC85111FDB96030148F0FC8";
   constant CPIX_NORMAL_INIT_00_BIT_02_C : bit_vector(255 downto 0) := x"47A0DA59A201983FCF7110A3F112FE12D7145035984D91F1D034A2BC94558440";
   constant CPIX_NORMAL_INIT_00_BIT_03_C : bit_vector(255 downto 0) := x"8C10558769867D524A5D71C0559A7D59630D69713A081B621254720500510440";
   constant CPIX_NORMAL_INIT_00_BIT_04_C : bit_vector(255 downto 0) := x"0F106C1842EF7512D09F2B8EFF2F6DFF73661F51837BE76F552097D704980E74";
   constant CPIX_NORMAL_INIT_00_BIT_05_C : bit_vector(255 downto 0) := x"07B014F615D3D5FEE048CA4EF041CEBB5F09099FC2B3C0BF322B9D8F57AB1B74";
   constant CPIX_NORMAL_INIT_00_BIT_06_C : bit_vector(255 downto 0) := x"0DE1242B24DBAC2BCD778ECBCE9706B36F474BF7A5BBB91D713DCFE246BD1E74";
   constant CPIX_NORMAL_INIT_00_BIT_07_C : bit_vector(255 downto 0) := x"28A15C6D7650B0A8F7C64DBEAD74BCED2F2650DED92FE4EE750BA7CF43DB1B74";
   constant CPIX_NORMAL_INIT_00_BIT_08_C : bit_vector(255 downto 0) := x"0321C0E82AECA6AF7B3F5B5E93188D59178E7ECF773392A21B7B559D370A5350";
   constant CPIX_NORMAL_INIT_00_BIT_09_C : bit_vector(255 downto 0) := x"1711E81D31AA439B128CFBFFEE8B1C6013E24F1B1AFFFB241D333FF4257C4650";
   constant CPIX_NORMAL_INIT_00_BIT_10_C : bit_vector(255 downto 0) := x"1380D77AEA68397E7C879BEA32A807C51B97F66769BF5E1839D56F3268756400";
   constant CPIX_NORMAL_INIT_00_BIT_11_C : bit_vector(255 downto 0) := x"1AB8A2C53B0E7054537BEDCE819D10393DD8734017EB8A066A501FB1703C4610";
   constant CPIX_NORMAL_INIT_00_BIT_12_C : bit_vector(255 downto 0) := x"11943D164D8F3A287212D833B70CAE0D09612B7651A5D2F224750C9D442A0710";
   constant CPIX_NORMAL_INIT_00_BIT_13_C : bit_vector(255 downto 0) := x"09D645DD70E415DD091B7CE0876F634C280A4C0A236C97526323569155180210";
   constant CPIX_NORMAL_INIT_00_BIT_14_C : bit_vector(255 downto 0) := x"43542BC470F02C1E76A4619376D4926A10784C635C4958970625222914560100";
   constant CPIX_NORMAL_INIT_01_BIT_00_C : bit_vector(255 downto 0) := x"DA45FFCF97D29EB2E0A3472FF71E47B9E981EF5C5DBA32B4ECC865649681F897";
   constant CPIX_NORMAL_INIT_01_BIT_01_C : bit_vector(255 downto 0) := x"55863F755814814E08DB81B95236213BFB69756850A94E8AD2D3BFF39993B885";
   constant CPIX_NORMAL_INIT_01_BIT_02_C : bit_vector(255 downto 0) := x"54429C40C7B507D7DF1C3907DE4492EBF5FC7ED0B1104D0EFB625354CB811565";
   constant CPIX_NORMAL_INIT_01_BIT_03_C : bit_vector(255 downto 0) := x"B5894254173BA06B6983843C7E632A48258F76A57C562010663783C54E8E319F";
   constant CPIX_NORMAL_INIT_01_BIT_04_C : bit_vector(255 downto 0) := x"10CE02554DB442803459A9AE7FF6425DA215D2FD4F8E45F8BBAA18B30886BDAE";
   constant CPIX_NORMAL_INIT_01_BIT_05_C : bit_vector(255 downto 0) := x"110A8F452764FF3C5767E75EF662BAF9AD4174C3A4C8E0ECEE40250FC48DD98F";
   constant CPIX_NORMAL_INIT_01_BIT_06_C : bit_vector(255 downto 0) := x"14C3E8025D601DCF1935F68E9CF04C8FA1B62F3BD5EDE1DBF5BDD33F7549881E";
   constant CPIX_NORMAL_INIT_01_BIT_07_C : bit_vector(255 downto 0) := x"08B0890333E539B26F3D36549B04DD84EE3FB47834B2DAA8DDF77B209A81ABE6";
   constant CPIX_NORMAL_INIT_01_BIT_08_C : bit_vector(255 downto 0) := x"051F5916F151BCC45888ADB59C29D9EA6B9F1BEE229F36A9D20A03D0D5873297";
   constant CPIX_NORMAL_INIT_01_BIT_09_C : bit_vector(255 downto 0) := x"472B4303A8C017A25A039DCD351BC69B561990B1FACAAEAFE8F9D5DA16842C41";
   constant CPIX_NORMAL_INIT_01_BIT_10_C : bit_vector(255 downto 0) := x"031EC110F32A2E98FD983C901FC23FE86AA5816F939FF9980F4D98D1410EA463";
   constant CPIX_NORMAL_INIT_01_BIT_11_C : bit_vector(255 downto 0) := x"02C98EC19D4CF0734EDB44AD7A457774220E3BDAECA2F1BD8113C6F707350AD3";
   constant CPIX_NORMAL_INIT_01_BIT_12_C : bit_vector(255 downto 0) := x"024787704EF7476934A394FA0BD90D802E5D5348A6950A4BDF3B54F0CDE845A2";
   constant CPIX_NORMAL_INIT_01_BIT_13_C : bit_vector(255 downto 0) := x"0596B66C7563A2B23B54B9711633F7A6009607CB2BA1B854807E2CBB385F61B0";
   constant CPIX_NORMAL_INIT_01_BIT_14_C : bit_vector(255 downto 0) := x"314B67654CDEB1756B45BB0109F103BC3A6C89652D53D65B2F2DE77493593D8D";
   constant CPIX_NORMAL_INIT_02_BIT_00_C : bit_vector(255 downto 0) := x"53393FBC5240984A8D196562E1B6619E425A5A3F83CDC69F6C923AED406B3884";
   constant CPIX_NORMAL_INIT_02_BIT_01_C : bit_vector(255 downto 0) := x"530DE9D086D84A2500E7025F3AB01BBC0FE802DBA3D8926A51EB030D3444064C";
   constant CPIX_NORMAL_INIT_02_BIT_02_C : bit_vector(255 downto 0) := x"43B5AFB2078A86C0E917CE8560EE81FC4A8B8C486B385B64268E1414D8A3B940";
   constant CPIX_NORMAL_INIT_02_BIT_03_C : bit_vector(255 downto 0) := x"B431D0BB4248FD322CB4372C5D101341CC386B6AC01D8122B0B910FA490786CD";
   constant CPIX_NORMAL_INIT_02_BIT_04_C : bit_vector(255 downto 0) := x"D54E02669A7DABF726BB91BD6427AEC1BACFCC8816D7FF5F04D1516C98E6DC9B";
   constant CPIX_NORMAL_INIT_02_BIT_05_C : bit_vector(255 downto 0) := x"81E775565E25F05BDC30E5D5AC15FCB5ECFD75545D3605AEE46414F3B093C0CB";
   constant CPIX_NORMAL_INIT_02_BIT_06_C : bit_vector(255 downto 0) := x"C5529E397CFB0FDEA226ACE2FC12F68ABB778EA6B74A0EEA2B36F4C3868442D9";
   constant CPIX_NORMAL_INIT_02_BIT_07_C : bit_vector(255 downto 0) := x"F5F95BAB9E352E900B719F5CA79C8DD5A3E2FA6F3A9A49508289C51399DFA81D";
   constant CPIX_NORMAL_INIT_02_BIT_08_C : bit_vector(255 downto 0) := x"609F92BA06DAECAD595C93AF0B7DCCD7B74905DC551BE641E767C02A5B59965F";
   constant CPIX_NORMAL_INIT_02_BIT_09_C : bit_vector(255 downto 0) := x"2A6942D78201CB16FE8DF59DC8EDD8BFECD0AB87F776B398522891750CE42567";
   constant CPIX_NORMAL_INIT_02_BIT_10_C : bit_vector(255 downto 0) := x"38D8C827C04738EAC20B87EBFF9696D004AE20F6C281B657210305AD8D21384F";
   constant CPIX_NORMAL_INIT_02_BIT_11_C : bit_vector(255 downto 0) := x"0C5944A80B8BE688BDE5DD5CAB06CBB6D107535BF529FE2A116A0B6640D8B70E";
   constant CPIX_NORMAL_INIT_02_BIT_12_C : bit_vector(255 downto 0) := x"58ED36E3371A7594DC6C9232159970CEA3AF0EDF3334EA11F4F6BDD065328D5C";
   constant CPIX_NORMAL_INIT_02_BIT_13_C : bit_vector(255 downto 0) := x"1411D769543AE19B4C8F9906DFD56724D5552EE949F19B9E1A8027FB3947CB40";
   constant CPIX_NORMAL_INIT_02_BIT_14_C : bit_vector(255 downto 0) := x"4F9C6CA4D583786309B7335BA629728A48FB18B6F86A3E70831A62D74BF780A6";
   constant CPIX_NORMAL_INIT_03_BIT_00_C : bit_vector(255 downto 0) := x"0D37CBC810545E106C915DA67C0671B217AE26E5DAC5A35014C5BD179BD4343C";
   constant CPIX_NORMAL_INIT_03_BIT_01_C : bit_vector(255 downto 0) := x"95ABA00FB414CBDCF1BEF13D47FFBEB1FCD02A80E078D77999265DC06C7C8419";
   constant CPIX_NORMAL_INIT_03_BIT_02_C : bit_vector(255 downto 0) := x"05217078D94B5522B37B9962C17EE722A7FE86AE1BC448FC85A47618C65EF70D";
   constant CPIX_NORMAL_INIT_03_BIT_03_C : bit_vector(255 downto 0) := x"E873D48277F81734077E0DDEDC012CD73993C45B84675FE719B1792A5C8C7C03";
   constant CPIX_NORMAL_INIT_03_BIT_04_C : bit_vector(255 downto 0) := x"4140F5E9401D436631A6D860304CC4194E3163C698D2D9E918A3EF7924092363";
   constant CPIX_NORMAL_INIT_03_BIT_05_C : bit_vector(255 downto 0) := x"411650C895EA5122597F6B61EBFA4FE5663A382EE97F76FC89252C5C8AD9AA56";
   constant CPIX_NORMAL_INIT_03_BIT_06_C : bit_vector(255 downto 0) := x"5065A00AAD81315D32F33C4156F2E4FE47970B32FB28C4FCE1ACBB4475E4C56B";
   constant CPIX_NORMAL_INIT_03_BIT_07_C : bit_vector(255 downto 0) := x"16D0DA15C487145E0B5BBC361F939E5C38AA5FF34F797365C1CF4430F2A394A5";
   constant CPIX_NORMAL_INIT_03_BIT_08_C : bit_vector(255 downto 0) := x"152613EB73864339EB0777579AF4B06023C4C1C589B7CE63D0A109D6A792AD99";
   constant CPIX_NORMAL_INIT_03_BIT_09_C : bit_vector(255 downto 0) := x"656F498E355A555F8DC0F041433ECC4C37C8004ED2A3E0E7492217CBA13CC6DE";
   constant CPIX_NORMAL_INIT_03_BIT_10_C : bit_vector(255 downto 0) := x"451A12FCA4435345EE4A1C9808EC9794FEF297905BE4875511BFF0180EBFB9D0";
   constant CPIX_NORMAL_INIT_03_BIT_11_C : bit_vector(255 downto 0) := x"514CF59280A8A406C2B360F4EF512B1E34E8F6DA217489B6799D75663A6F7B61";
   constant CPIX_NORMAL_INIT_03_BIT_12_C : bit_vector(255 downto 0) := x"5009242A847F6F5460FDFA2A257E7CD64E21894F8660BFDD478FF28741F2D544";
   constant CPIX_NORMAL_INIT_03_BIT_13_C : bit_vector(255 downto 0) := x"1076833DCA387CF47E66390E9909DB190BCF27208A926F5642780E4BEF2EC938";
   constant CPIX_NORMAL_INIT_03_BIT_14_C : bit_vector(255 downto 0) := x"1E03618F7D6A383321E4A2FD9A436B736D8A65268ECF011745C3FB52141B8EE0";
   constant CPIX_NORMAL_INIT_04_BIT_00_C : bit_vector(255 downto 0) := x"9EF3CD229D72A4106FB54B085AD22D04965A3DF7B53747089BBF8321A03F2A8E";
   constant CPIX_NORMAL_INIT_04_BIT_01_C : bit_vector(255 downto 0) := x"75F3DA1837C1E9244D4546266234AA765EF62E960FC2F8103A2459EB4AACF5C5";
   constant CPIX_NORMAL_INIT_04_BIT_02_C : bit_vector(255 downto 0) := x"7081A44F95E9621FE884AA50A7C729AD297814B4576942C2A3D4ED1B9BD26164";
   constant CPIX_NORMAL_INIT_04_BIT_03_C : bit_vector(255 downto 0) := x"A5AD0A056DDE281DA14F1632915F4959CE541F9A4254AEA92592452BC06CB5F2";
   constant CPIX_NORMAL_INIT_04_BIT_04_C : bit_vector(255 downto 0) := x"8E9CB13AA0B4C141463DE6FAAEFA27AA4465671632527DF5D790FD2CB6A193DA";
   constant CPIX_NORMAL_INIT_04_BIT_05_C : bit_vector(255 downto 0) := x"ACE5BF377B6263F436F25E28552388FDA864F9740721AA5EDA51D35AE045B19B";
   constant CPIX_NORMAL_INIT_04_BIT_06_C : bit_vector(255 downto 0) := x"CACE7FEFD4FCC8799F2B618C01E8FCCC1CDE1A2DEA70B10B807CC461355CF682";
   constant CPIX_NORMAL_INIT_04_BIT_07_C : bit_vector(255 downto 0) := x"D85FAD18AEDC3CAE5BD9D3DD30C27250D10DD097B132165BD397F6BF99C557E6";
   constant CPIX_NORMAL_INIT_04_BIT_08_C : bit_vector(255 downto 0) := x"DA3F75971523F6A56236569EF83C7516AC6B6C2EB0445DD9329B66D7D22D73BF";
   constant CPIX_NORMAL_INIT_04_BIT_09_C : bit_vector(255 downto 0) := x"EDB5E654989AC46BFF3B6E7CCB1FC395631D0CD493076A6744A4B8644C263D6E";
   constant CPIX_NORMAL_INIT_04_BIT_10_C : bit_vector(255 downto 0) := x"017198FD4810EF6DA55C85529F39673B4C42111A442298E2D4A64C120E9074BA";
   constant CPIX_NORMAL_INIT_04_BIT_11_C : bit_vector(255 downto 0) := x"B657053F671E63DAAE334DD7FEAD58D80706798D418A3D296044A3908B2E50ED";
   constant CPIX_NORMAL_INIT_04_BIT_12_C : bit_vector(255 downto 0) := x"885EC9FB14EDB6EF4E5B0E30BDCC0713FF31AB698AE3B2406D674A5880F622B4";
   constant CPIX_NORMAL_INIT_04_BIT_13_C : bit_vector(255 downto 0) := x"E366623618EDA8D63596EB57838ED7B956C985145C7FEECE1ED7756FB0DB7141";
   constant CPIX_NORMAL_INIT_04_BIT_14_C : bit_vector(255 downto 0) := x"25C4EBDF0690DE2CFEC4388D4BE83B50914A07DC3C0DA26B359FBE2FD144897D";
   constant CPIX_NORMAL_INIT_05_BIT_00_C : bit_vector(255 downto 0) := x"8DF4E16DB415340F9DF7DAFF3D3EDB667A1CB86CD298C3A347B86093C2F87D53";
   constant CPIX_NORMAL_INIT_05_BIT_01_C : bit_vector(255 downto 0) := x"15454E75B6392DB4E2719795F71978EAD5A2AABD287F1EF3B28B417C6BCC4808";
   constant CPIX_NORMAL_INIT_05_BIT_02_C : bit_vector(255 downto 0) := x"47519BF085380D1D0433E4C891BCB450AC974629E1E9F16E740576ACD5152C14";
   constant CPIX_NORMAL_INIT_05_BIT_03_C : bit_vector(255 downto 0) := x"BE6F0E55EAD719CE75417581EBE25F0C19A4CE230F7F08F46BB7DE14464CE7B2";
   constant CPIX_NORMAL_INIT_05_BIT_04_C : bit_vector(255 downto 0) := x"F32235BE404CFF3C97846EB39C9FAF6A1D39CEDBC3539FA66964092FC8EEA046";
   constant CPIX_NORMAL_INIT_05_BIT_05_C : bit_vector(255 downto 0) := x"D553E93B2A67773C27E51C76BB0433DFE2E50B14B873E636DCF40222AAF59E37";
   constant CPIX_NORMAL_INIT_05_BIT_06_C : bit_vector(255 downto 0) := x"F172630D86B94BC32FECEECA00AAE2F88D5D1C7D99B0BC19EFE5131DFF3984D9";
   constant CPIX_NORMAL_INIT_05_BIT_07_C : bit_vector(255 downto 0) := x"FB36FBC227DA8D8A93A80B261DEDD241058F6A53D7EE63E09C3A86F184E7B726";
   constant CPIX_NORMAL_INIT_05_BIT_08_C : bit_vector(255 downto 0) := x"2C5082EEC3598FDD1169A69CE8B0CCF266C667A0D60AC8AE558B3AA2A4A4E33E";
   constant CPIX_NORMAL_INIT_05_BIT_09_C : bit_vector(255 downto 0) := x"598D79C73409F37ED00C1056B08A563DBFED94B3AE7397E2E0D5ECE6E3C18FAE";
   constant CPIX_NORMAL_INIT_05_BIT_10_C : bit_vector(255 downto 0) := x"4E84E3D0B1854C7EE554653B4A80F89CF10D44CFD43AED9AEBFA826DC77CF605";
   constant CPIX_NORMAL_INIT_05_BIT_11_C : bit_vector(255 downto 0) := x"54B567C26065899115CB85CFED7D81918AF3E963E3A366B5D9DB056DF4DA8E38";
   constant CPIX_NORMAL_INIT_05_BIT_12_C : bit_vector(255 downto 0) := x"2280E9A71E7DAD5F4A7F42882F779621B7B46DA1820D4A5D1326D3972B00E1FD";
   constant CPIX_NORMAL_INIT_05_BIT_13_C : bit_vector(255 downto 0) := x"46215753F63B7C8232315AC9B917C2DB21E5D4BAD6864168E6FFB767796E5D70";
   constant CPIX_NORMAL_INIT_05_BIT_14_C : bit_vector(255 downto 0) := x"74FE87A129F48C75B623904F7F906D1F15C29A6E5E1B729F98294C936F19D098";
   constant CPIX_NORMAL_INIT_06_BIT_00_C : bit_vector(255 downto 0) := x"E9846646F29616894C325ADC27F4CCBEE99E1ECD654CB9806C711DCBE5DEF51E";
   constant CPIX_NORMAL_INIT_06_BIT_01_C : bit_vector(255 downto 0) := x"F89E7BBD01E42C324B9C8BB23B7509C6D1E2FD4FA915B63FBF3BCC90DE515D76";
   constant CPIX_NORMAL_INIT_06_BIT_02_C : bit_vector(255 downto 0) := x"CE1F6BAC8D645CE9A28AC564E4DFDDE4D7628C517DCA4295F1B944D9FB5E1367";
   constant CPIX_NORMAL_INIT_06_BIT_03_C : bit_vector(255 downto 0) := x"0AA6560EF128A39BD5604C2F27EB9A7E02978F7379E71D9833E0F7D56B9411CF";
   constant CPIX_NORMAL_INIT_06_BIT_04_C : bit_vector(255 downto 0) := x"21ECCA57294AF47C86D5C359A2D6D8C607D09D5BAAAB2BD30C7441B24C7B3C0E";
   constant CPIX_NORMAL_INIT_06_BIT_05_C : bit_vector(255 downto 0) := x"386D4FDD1F9549EDED874AEE2A6C8BB081D359674DF432A081CDA296DCCC377C";
   constant CPIX_NORMAL_INIT_06_BIT_06_C : bit_vector(255 downto 0) := x"256E837F51DB4A18FBCB78D1A125CFF0B9569DA0DEDA70646F72E865A176389A";
   constant CPIX_NORMAL_INIT_06_BIT_07_C : bit_vector(255 downto 0) := x"1BC5CD9C22BAAE5B60BA2E826E5A0976A453E1BB34244A54FB19884B92309877";
   constant CPIX_NORMAL_INIT_06_BIT_08_C : bit_vector(255 downto 0) := x"1C4FB125E003F122C0838E7FA1EC1C5AB20488170483B67DD87AC60D98B29382";
   constant CPIX_NORMAL_INIT_06_BIT_09_C : bit_vector(255 downto 0) := x"1B6EA4C1051070E8B75CCD1FBD50C82A20C60C58177AB59ACD171AF5E52DF6A9";
   constant CPIX_NORMAL_INIT_06_BIT_10_C : bit_vector(255 downto 0) := x"BFBDAF48C72E865437CFF860847B176306139AEBFF1056C014ADDFFF8FC7F254";
   constant CPIX_NORMAL_INIT_06_BIT_11_C : bit_vector(255 downto 0) := x"0E20ADD1FE68F6DD4C122B708583FA786F86C3E67F6638384FD96DFA2FCE3C42";
   constant CPIX_NORMAL_INIT_06_BIT_12_C : bit_vector(255 downto 0) := x"60E90C02949761AFD46C6954CEBBB2B3642E91FABA4DD12F3503AB19B7272571";
   constant CPIX_NORMAL_INIT_06_BIT_13_C : bit_vector(255 downto 0) := x"108AB4EE5C7B5910C4CC965C7CAE372D60097B8051F964DEBDFB0CFDB5974E80";
   constant CPIX_NORMAL_INIT_06_BIT_14_C : bit_vector(255 downto 0) := x"39F691D968234C3DC4EDF0AB5402567B7073A00EFE9B320D1631178E95EDB815";
   constant CPIX_NORMAL_INIT_07_BIT_00_C : bit_vector(255 downto 0) := x"EE49F5C11F714F2FBDBAD9DE8D52A9FB861E3CEC984D6396C04EAFD3C4F874E7";
   constant CPIX_NORMAL_INIT_07_BIT_01_C : bit_vector(255 downto 0) := x"D2C1C7E42DDEB07ED96031448376F5F5C6F75CAA8CE4D78E0ACAEED6B5AE504E";
   constant CPIX_NORMAL_INIT_07_BIT_02_C : bit_vector(255 downto 0) := x"44051558FF452F45A5D326AB07FB1E49A25EB9CEB195646994362AD5A73BD25C";
   constant CPIX_NORMAL_INIT_07_BIT_03_C : bit_vector(255 downto 0) := x"BCA7735DA660C09D692BFA90736E4F30583A3CEC53A4FBBC97E4406A44B4FF7F";
   constant CPIX_NORMAL_INIT_07_BIT_04_C : bit_vector(255 downto 0) := x"31533953FF73FD92731412B3315E69790E07DF6DB7C22C153B4571B0ED7547C6";
   constant CPIX_NORMAL_INIT_07_BIT_05_C : bit_vector(255 downto 0) := x"3447077C3201B1908226F8C97747595C32927FAB6CCB6D07FD8FEEDD75AFF972";
   constant CPIX_NORMAL_INIT_07_BIT_06_C : bit_vector(255 downto 0) := x"76517976CC4114D9CDE784524B4237A20E4CFA0A0BB421572328BA0DAD21BFF9";
   constant CPIX_NORMAL_INIT_07_BIT_07_C : bit_vector(255 downto 0) := x"172DE240B7895772A175953B173467ED008E638ECEF05A2957EED20F96F832F0";
   constant CPIX_NORMAL_INIT_07_BIT_08_C : bit_vector(255 downto 0) := x"0733586D435EB9CF3A0E853D754F5A93A99B106F2A3F736FD6D8EB208F052D10";
   constant CPIX_NORMAL_INIT_07_BIT_09_C : bit_vector(255 downto 0) := x"2D2768BA70D7C5E84E636389622663BF85A6B514BF103442615B4EFCE1E134F1";
   constant CPIX_NORMAL_INIT_07_BIT_10_C : bit_vector(255 downto 0) := x"3463028D1648AEE18920741E360F3527A8B930CC17F0C6D54190FCB0836B8360";
   constant CPIX_NORMAL_INIT_07_BIT_11_C : bit_vector(255 downto 0) := x"221334F5FA76970C9015DD808975452CA41CDA0A2C00BE31A8AA621749DF06E9";
   constant CPIX_NORMAL_INIT_07_BIT_12_C : bit_vector(255 downto 0) := x"2745018359350DD9D1646FFE29FE76303D01AEF7BF8D4D980C733BAD3FF4A22D";
   constant CPIX_NORMAL_INIT_07_BIT_13_C : bit_vector(255 downto 0) := x"07102A3D811B1AA7A0990AC07BF1EA357FBD6C7D1EC301E996C31582E39E07D2";
   constant CPIX_NORMAL_INIT_07_BIT_14_C : bit_vector(255 downto 0) := x"07BD100A6C5795AB7AB33C9D1BD41B1E4947ED71DC59AFA6C69D304A38CE7F1F";
   constant CPIX_NORMAL_INIT_08_BIT_00_C : bit_vector(255 downto 0) := x"7DC7D837F10D45C0718CA4D1DBD1EA6E6C6134553FE1A2E837AFF045F2332E16";
   constant CPIX_NORMAL_INIT_08_BIT_01_C : bit_vector(255 downto 0) := x"E491D9E1435B28168FD8EE679BBA42819D53C2DBA798E09DAD9C831AE2EF349A";
   constant CPIX_NORMAL_INIT_08_BIT_02_C : bit_vector(255 downto 0) := x"0AEF19994A855D59365829DB544CA5499E96EE54BCE15F9D83DAFFE83012A805";
   constant CPIX_NORMAL_INIT_08_BIT_03_C : bit_vector(255 downto 0) := x"A4FC016012CF54BC352F3625E8A898D2586F8769216559DCF14528E49273FF39";
   constant CPIX_NORMAL_INIT_08_BIT_04_C : bit_vector(255 downto 0) := x"21310A237D0ED5795B4D374C3BA3BF33E66A9701FAF119A3CF788C579A5FB2CD";
   constant CPIX_NORMAL_INIT_08_BIT_05_C : bit_vector(255 downto 0) := x"99C00971BAF72871452A48579C9C22BDB7C92653B74877CDF91071268B53D28E";
   constant CPIX_NORMAL_INIT_08_BIT_06_C : bit_vector(255 downto 0) := x"42B497AD46891AA3ECD83F44CB56559AD1452AF1A03678531F2663A4BE3C8019";
   constant CPIX_NORMAL_INIT_08_BIT_07_C : bit_vector(255 downto 0) := x"A60731E2B355936E8A165F0D1329778BB61F822BEB298FFFD6D3E462376EF969";
   constant CPIX_NORMAL_INIT_08_BIT_08_C : bit_vector(255 downto 0) := x"DDA06CDA78B45DE9CE51253133E3B3D25B58D39B282CF73BE7084CA37B5B8EFF";
   constant CPIX_NORMAL_INIT_08_BIT_09_C : bit_vector(255 downto 0) := x"281A42B210B4F761965A557A6DD93D6A20719835DFD0282534A40D3C1EE62DBC";
   constant CPIX_NORMAL_INIT_08_BIT_10_C : bit_vector(255 downto 0) := x"34F075185756169935341D1D83D4FD0DA7648D7D21A1425955ED93112F34DED8";
   constant CPIX_NORMAL_INIT_08_BIT_11_C : bit_vector(255 downto 0) := x"056F402C6FD7D0E67013D5DD4EA21DC37C503131880A8351C0CF0CF93350B9E6";
   constant CPIX_NORMAL_INIT_08_BIT_12_C : bit_vector(255 downto 0) := x"AFBE0E52DD8F7896C1D8AD1BCE09311529A6297A218C32908515FF2C0C4CDE30";
   constant CPIX_NORMAL_INIT_08_BIT_13_C : bit_vector(255 downto 0) := x"3779A193D173122167B06EEEA8ACB1E912ACF76A7E6729AF9F00E69A6F123416";
   constant CPIX_NORMAL_INIT_08_BIT_14_C : bit_vector(255 downto 0) := x"8646609D543AF6E41FE500E78C18399E5F27C7BF8EF91DAEB206357094932BB2";
   constant CPIX_NORMAL_INIT_09_BIT_00_C : bit_vector(255 downto 0) := x"7D0210A44E5CB2E73C5881F777DFB9FBD25174DD8A71FF6FC8370CE7E348FECA";
   constant CPIX_NORMAL_INIT_09_BIT_01_C : bit_vector(255 downto 0) := x"B9DB0010477E1FDDDCD88F0E75F31E601C18EB4551A758F95AD5AC2DD13E2E0C";
   constant CPIX_NORMAL_INIT_09_BIT_02_C : bit_vector(255 downto 0) := x"7C606A4938B165FE9000CC96B54917EEDC23C157BD943311AC77E37A10069896";
   constant CPIX_NORMAL_INIT_09_BIT_03_C : bit_vector(255 downto 0) := x"9A760CF094C851767AD096AC009446F2F89235CA17750A1D831F37FF2D5667B7";
   constant CPIX_NORMAL_INIT_09_BIT_04_C : bit_vector(255 downto 0) := x"81BC57F39A025EDD9D32AF71F903711334384A87F970AE8999B9EBCC5CFED999";
   constant CPIX_NORMAL_INIT_09_BIT_05_C : bit_vector(255 downto 0) := x"D8F529228BFF5E6F3B9B3858285EEA315A3CAE7C23E41C8133331D5F8481EFA3";
   constant CPIX_NORMAL_INIT_09_BIT_06_C : bit_vector(255 downto 0) := x"B58D75A82FAEECBFF620AEF5F4C17A9787FB1CCB681E91B10503FCC0BAB1E4E5";
   constant CPIX_NORMAL_INIT_09_BIT_07_C : bit_vector(255 downto 0) := x"E2D4E2BB88F613908DADA7F01BE4DCEC239FA3D2F74EA3E71B51A0092B0C7745";
   constant CPIX_NORMAL_INIT_09_BIT_08_C : bit_vector(255 downto 0) := x"A28C4AAE7A72936A42364D4FBB289D37795D1F69777DC2A8EAC00FF53B235238";
   constant CPIX_NORMAL_INIT_09_BIT_09_C : bit_vector(255 downto 0) := x"ECA2DA76B8792270D6D09789A0653D9ABEAA1B9A68BC3BF1B4CF07BEA01F9727";
   constant CPIX_NORMAL_INIT_09_BIT_10_C : bit_vector(255 downto 0) := x"55472B538785EBE365D00644BCAF79F2DD2737F48036375887FB1AD3287F0BDA";
   constant CPIX_NORMAL_INIT_09_BIT_11_C : bit_vector(255 downto 0) := x"8E6D332B05770FFF7D6B16A9395EE6CCDCFC4F0B74E2E32FEFECC9F27691A2D4";
   constant CPIX_NORMAL_INIT_09_BIT_12_C : bit_vector(255 downto 0) := x"908477FDE182ABDF5335FCF2DF7CACBE61E862CB45A94E459FF2A5F0046B521B";
   constant CPIX_NORMAL_INIT_09_BIT_13_C : bit_vector(255 downto 0) := x"BC5F6D3C385D4E385784E8E289C1E6291F738728B98E663F944BD1B8E76ACF82";
   constant CPIX_NORMAL_INIT_09_BIT_14_C : bit_vector(255 downto 0) := x"5C73E531ACCEE3FB112CD755A3FD09F1AAECE5640EC5D1B331DEEC910A8B6310";
   constant CPIX_NORMAL_INIT_0A_BIT_00_C : bit_vector(255 downto 0) := x"9532A91A717AC35B0DE63D7E4AF066E19A90757BC6BF39E40FA2403B814DDCE4";
   constant CPIX_NORMAL_INIT_0A_BIT_01_C : bit_vector(255 downto 0) := x"98EEDAA9530CA753BB9CBC7AF2F26604EF365F0E1D47EDEFCDC25F655E23728A";
   constant CPIX_NORMAL_INIT_0A_BIT_02_C : bit_vector(255 downto 0) := x"BAF0D76FEDAD5563AD17FF17BE4EA5F32F6980A31F2DCEE0C67EF6A268244371";
   constant CPIX_NORMAL_INIT_0A_BIT_03_C : bit_vector(255 downto 0) := x"07978970E1F850DA11BE7E3A5185B72D7C9BDB6AD6FC5225542D74F0BCFBCA0D";
   constant CPIX_NORMAL_INIT_0A_BIT_04_C : bit_vector(255 downto 0) := x"43A74ED2E1A8FEDAE40F76DF96AFD4396986396425D60CBE9594F8FC8805756D";
   constant CPIX_NORMAL_INIT_0A_BIT_05_C : bit_vector(255 downto 0) := x"A81DB827148B4334DA916B5AA968076DE7E1FF70401C1919E8D9BF3297E81A6A";
   constant CPIX_NORMAL_INIT_0A_BIT_06_C : bit_vector(255 downto 0) := x"C5B763B353E03BA3D3D29F55DBA55B92E8ABF877424E06F6EAEA1A92C434E2D7";
   constant CPIX_NORMAL_INIT_0A_BIT_07_C : bit_vector(255 downto 0) := x"0533D4AA28C8375BF37FBCAD790BFC4083E40F89C078AA42D020BC7BCB2F5D79";
   constant CPIX_NORMAL_INIT_0A_BIT_08_C : bit_vector(255 downto 0) := x"686DA17C393BCC10E63C118DE0C099BD2636858B1ACCDC1CC8748824AC5B5BAD";
   constant CPIX_NORMAL_INIT_0A_BIT_09_C : bit_vector(255 downto 0) := x"CFFABCA78374DE0EC8BC3B4A867AB919ED14F633FCF5BC3DF90FE112D1BE8CF9";
   constant CPIX_NORMAL_INIT_0A_BIT_10_C : bit_vector(255 downto 0) := x"AF5341F36424B1EEF6315ADCE8F39398EC8BAF9C811979B6F53B7FB1AF281537";
   constant CPIX_NORMAL_INIT_0A_BIT_11_C : bit_vector(255 downto 0) := x"D48CFA4BE9967C1BEC4E980B6D6C9E62F2C7B39A406239E7BF21B3CDC1FC5ED4";
   constant CPIX_NORMAL_INIT_0A_BIT_12_C : bit_vector(255 downto 0) := x"9F7ACE3578B3CD12915851E6619932F2075A4C69A24B937A1D8F0141B947FAF3";
   constant CPIX_NORMAL_INIT_0A_BIT_13_C : bit_vector(255 downto 0) := x"4C07B932F660CF89F668917874426D85B968FAEA9F2F686E3BD739B873F32E05";
   constant CPIX_NORMAL_INIT_0A_BIT_14_C : bit_vector(255 downto 0) := x"0326A14D82CC69AD66E9438A6B1DC6EED695198731E5C21F6CBB1786F75196D1";
   constant CPIX_NORMAL_INIT_0B_BIT_00_C : bit_vector(255 downto 0) := x"6A0C55DE17FDD658218FECC9A48EFF05781805C14C620100F548F1174C708283";
   constant CPIX_NORMAL_INIT_0B_BIT_01_C : bit_vector(255 downto 0) := x"D2D58F5688FF06D4104C59B552C29E8A7FAFD12C61B33989B5D8486A8C5BC0F5";
   constant CPIX_NORMAL_INIT_0B_BIT_02_C : bit_vector(255 downto 0) := x"701C5733E78E82325F474C9308C357C6D434654D3F2822F28C359871FDE15E49";
   constant CPIX_NORMAL_INIT_0B_BIT_03_C : bit_vector(255 downto 0) := x"8B8F08AA44BC4E7329A8E46A13B3B1DC2F767E40FE365053EED8FFC975FB34F1";
   constant CPIX_NORMAL_INIT_0B_BIT_04_C : bit_vector(255 downto 0) := x"AE6F38581B66EBE8F01033B1BBEE1E80837ED4626DB80F0F83A293AB8EEF7D9D";
   constant CPIX_NORMAL_INIT_0B_BIT_05_C : bit_vector(255 downto 0) := x"E763361EAC971FDA4CDD3D3B2A6E5BD54D3EED3652B4AA6DCA9A00605A0FA3EA";
   constant CPIX_NORMAL_INIT_0B_BIT_06_C : bit_vector(255 downto 0) := x"BF127A593C1B04B7D478DB9260CFE03E5CBBF8E1A8FDB08940448DDCA819AF91";
   constant CPIX_NORMAL_INIT_0B_BIT_07_C : bit_vector(255 downto 0) := x"BECB0A29EFCBE51D187EE28CD1A785C8C24BCCC044DB586812B6B8A2B3096113";
   constant CPIX_NORMAL_INIT_0B_BIT_08_C : bit_vector(255 downto 0) := x"1DA17204851CECADF54E769390FBE3A2421678C2882992F1E885CF51E0A1FB5D";
   constant CPIX_NORMAL_INIT_0B_BIT_09_C : bit_vector(255 downto 0) := x"33C380E26E87B56F0A3550C7BA4F6BF8A25114E1075533789E00C0D933284BF2";
   constant CPIX_NORMAL_INIT_0B_BIT_10_C : bit_vector(255 downto 0) := x"65BC8124F84AF654CF47D02264E43EFDE967227578735EDB258D9505EAD5C6B5";
   constant CPIX_NORMAL_INIT_0B_BIT_11_C : bit_vector(255 downto 0) := x"23759B72393BB1196C506C3284D383534773E58B8022B1EFE8F32EA294029302";
   constant CPIX_NORMAL_INIT_0B_BIT_12_C : bit_vector(255 downto 0) := x"1D589441ACD78D2A03BC2BB389B272BA74D83BBA605D95C118AE6A2B82284853";
   constant CPIX_NORMAL_INIT_0B_BIT_13_C : bit_vector(255 downto 0) := x"20785843772B621FEA6C1ACF7FE190195A190B537799B083CB93466AA108E38A";
   constant CPIX_NORMAL_INIT_0B_BIT_14_C : bit_vector(255 downto 0) := x"2A64EAFCC16E9C4619C2FF3495E53B269B6C584ED70065BF6EFB93456DF717FE";
   constant CPIX_NORMAL_INIT_0C_BIT_00_C : bit_vector(255 downto 0) := x"436C3C07E8574F5CC2889E1B253C3EFA934F90ECA8590F7106C80D1345DDA843";
   constant CPIX_NORMAL_INIT_0C_BIT_01_C : bit_vector(255 downto 0) := x"0BC16EE4BD0F8448F4F5279344AE8BAEA30A619DA35677DF4BCBD5FF9C9428D4";
   constant CPIX_NORMAL_INIT_0C_BIT_02_C : bit_vector(255 downto 0) := x"173CED05D64446F467E4E0E9BF5CC222F2F3848130D166920EEB11B870292F16";
   constant CPIX_NORMAL_INIT_0C_BIT_03_C : bit_vector(255 downto 0) := x"A45AC272C50F4E087394E87F42A3D3C5165BF343FF5E2273CDDBB0710105F0C6";
   constant CPIX_NORMAL_INIT_0C_BIT_04_C : bit_vector(255 downto 0) := x"103BA20DC746479CC5DAC9CF4C9EB35B49F0737535660B1941E0288A09B354D5";
   constant CPIX_NORMAL_INIT_0C_BIT_05_C : bit_vector(255 downto 0) := x"C403F74F7332582D3DA7FF744B0C8800C056FCA3D809032D97A5A2B4487F7F8D";
   constant CPIX_NORMAL_INIT_0C_BIT_06_C : bit_vector(255 downto 0) := x"CB9366388322BD57F3ACE3983B1568757CEB2A09F881F862E9066B6959D4D7F9";
   constant CPIX_NORMAL_INIT_0C_BIT_07_C : bit_vector(255 downto 0) := x"9D74261FA996DF9B0A704D65358C7375AA9E5696D480248BD71C5F40D4D02E7A";
   constant CPIX_NORMAL_INIT_0C_BIT_08_C : bit_vector(255 downto 0) := x"CE4C5570C490173F1071D40F8F7D7FA6F6C43AD8F02904A293848F48814E910D";
   constant CPIX_NORMAL_INIT_0C_BIT_09_C : bit_vector(255 downto 0) := x"1911B02C10F17791062B3B8D9A2397D8E4F3122E569CAA37AC774CA3E82D9993";
   constant CPIX_NORMAL_INIT_0C_BIT_10_C : bit_vector(255 downto 0) := x"446D430F87CCFDDFEFFE1244326CE110536189E2A2EBFAEBD4FFA53FE9193220";
   constant CPIX_NORMAL_INIT_0C_BIT_11_C : bit_vector(255 downto 0) := x"3CBE9179E00FF93D2BBE2D780BD50F9071FEB38239B2EFD80CFFB1F818A4650C";
   constant CPIX_NORMAL_INIT_0C_BIT_12_C : bit_vector(255 downto 0) := x"297159ADD647BAD99B9D64E6E3534CEE5E73054BC88A17D38F7B587A5E736F53";
   constant CPIX_NORMAL_INIT_0C_BIT_13_C : bit_vector(255 downto 0) := x"6C4401D26BCED0402303EFD63D35E3EC8EE7EF9E54F4ABA78E73C62E21F8D011";
   constant CPIX_NORMAL_INIT_0C_BIT_14_C : bit_vector(255 downto 0) := x"3B117F1B9C0050F8ABF897DB5A5C01B3122D1F47172BC4FDC637BDE6CFD04637";
   constant CPIX_NORMAL_INIT_0D_BIT_00_C : bit_vector(255 downto 0) := x"53697ADAD796DFC304E22987E9863B688F0FE4B2CC734D0AF694159B0F0F7452";
   constant CPIX_NORMAL_INIT_0D_BIT_01_C : bit_vector(255 downto 0) := x"465252DC46E2AB8BAF0E2A485E889ECB407FDDFDE24638AD12B1C046B5263B81";
   constant CPIX_NORMAL_INIT_0D_BIT_02_C : bit_vector(255 downto 0) := x"5878829F55869885C5E7B8006695FDC2ACD8D39CB0BFFB21F53A8D8BB636680C";
   constant CPIX_NORMAL_INIT_0D_BIT_03_C : bit_vector(255 downto 0) := x"A009DD5C4F74549CFE4348F48D7F86CEA2227C1024F008FB543F8ABB9608EECC";
   constant CPIX_NORMAL_INIT_0D_BIT_04_C : bit_vector(255 downto 0) := x"0DC3F8D594D4364F5C8635D9FE243FF1902DE232E11B2787D54D8669F711B50D";
   constant CPIX_NORMAL_INIT_0D_BIT_05_C : bit_vector(255 downto 0) := x"5E852CC714E6F69217BF82323582ADA6FDA2953F3589BCA900890CF0D05ADB35";
   constant CPIX_NORMAL_INIT_0D_BIT_06_C : bit_vector(255 downto 0) := x"0863789DE1132EDE6617B7CA31DC4690BE8FA08B6AD1E61394063C23E02ABA41";
   constant CPIX_NORMAL_INIT_0D_BIT_07_C : bit_vector(255 downto 0) := x"138AE053F4BE92914918CA89DCB9379E69059EC94CB9944964A872C840167A68";
   constant CPIX_NORMAL_INIT_0D_BIT_08_C : bit_vector(255 downto 0) := x"02E030DBDB535852FC45404AAE460D09F401840A91BD3FBA8407F9B4423526DC";
   constant CPIX_NORMAL_INIT_0D_BIT_09_C : bit_vector(255 downto 0) := x"039A68C9C925F567017642542F51E980DB6A26E1F0F353BBC6B67654A0044899";
   constant CPIX_NORMAL_INIT_0D_BIT_10_C : bit_vector(255 downto 0) := x"CEBEDAD6C9FE35D0A17A1DF9906977640E3FF1EBAB94384488753BCF57BF294E";
   constant CPIX_NORMAL_INIT_0D_BIT_11_C : bit_vector(255 downto 0) := x"45E8192098A7E706FFE87985BF68B7B370B1531D099A3F55C572955BFFDD3F95";
   constant CPIX_NORMAL_INIT_0D_BIT_12_C : bit_vector(255 downto 0) := x"7945FDC240E015599264976F684799FBF27029B16D836660F1F89B9BDF499F4F";
   constant CPIX_NORMAL_INIT_0D_BIT_13_C : bit_vector(255 downto 0) := x"5605D5898F70FDBD66F16F9B22821211A424B5F1976D76E52FB589B95F6F19E6";
   constant CPIX_NORMAL_INIT_0D_BIT_14_C : bit_vector(255 downto 0) := x"0AC7BE7C8202F3D629C01D5F25F44EA2E531ADA7FF0198DF3631054D773D6BCE";
   constant CPIX_NORMAL_INIT_0E_BIT_00_C : bit_vector(255 downto 0) := x"3FD7BD47E10B125B3D3BCA5DC6A16D924AEF8B57330558E14BCB146A91CA1290";
   constant CPIX_NORMAL_INIT_0E_BIT_01_C : bit_vector(255 downto 0) := x"3104FCC76C0030395364CD878B2517D1F0999425745640766A5226290D31D883";
   constant CPIX_NORMAL_INIT_0E_BIT_02_C : bit_vector(255 downto 0) := x"58603181987768784A93B313583BACFEC3243BF0D571016F0C4A924B904D47C8";
   constant CPIX_NORMAL_INIT_0E_BIT_03_C : bit_vector(255 downto 0) := x"E7C90DE108257865B64E8805CA8FCBA4936FB838399C9F8DB01186A088BB1FCE";
   constant CPIX_NORMAL_INIT_0E_BIT_04_C : bit_vector(255 downto 0) := x"44E80336A13BA8339F7AA42D79F016664F8E60767B17AE54AC872627172B9408";
   constant CPIX_NORMAL_INIT_0E_BIT_05_C : bit_vector(255 downto 0) := x"0A4D8240282A885E78F5A4DF29B2107FEBE294EEBDFCB7B62E02C5AA8BD65F7C";
   constant CPIX_NORMAL_INIT_0E_BIT_06_C : bit_vector(255 downto 0) := x"14F961FCA91C115D04DA9A215D43766E1D1B0DD09B8904E79C825106EFFBDE86";
   constant CPIX_NORMAL_INIT_0E_BIT_07_C : bit_vector(255 downto 0) := x"4514C0FD7E9A9129E0FCEA40678D1986766EF8EDB74800EF860CE6915A0CCA14";
   constant CPIX_NORMAL_INIT_0E_BIT_08_C : bit_vector(255 downto 0) := x"CC97D29F57516C7A588C1BEB2B1A6CBEF338B290AD8F5814D1CE493619E22701";
   constant CPIX_NORMAL_INIT_0E_BIT_09_C : bit_vector(255 downto 0) := x"C473DD3D8E6643E4CEFA06545E24244D391662CE70E8FFF4ED63A8565E30EA12";
   constant CPIX_NORMAL_INIT_0E_BIT_10_C : bit_vector(255 downto 0) := x"88809AD61E54B4A4472FBE44E16DB36660168741EAB0DF51915F68DB845E6811";
   constant CPIX_NORMAL_INIT_0E_BIT_11_C : bit_vector(255 downto 0) := x"8C3157B1A68804884CE145448FA90F138D91CDDD3D1C422B35D3F6FB0179ADC7";
   constant CPIX_NORMAL_INIT_0E_BIT_12_C : bit_vector(255 downto 0) := x"4BF744438DB9EA7EDFEB91B334B2C38540E07B4A0B8BDCB60FFBAE34DC4D4DA3";
   constant CPIX_NORMAL_INIT_0E_BIT_13_C : bit_vector(255 downto 0) := x"7EEFCEB63CB16EB306FCA14E0053B982933DA54B4663954DAD4BC7B8153BF258";
   constant CPIX_NORMAL_INIT_0E_BIT_14_C : bit_vector(255 downto 0) := x"60D3352EB9A66B13E6B12682C9ABC82CF47CC3A34F0135881BC4F4BC2EAE52EA";
   constant CPIX_NORMAL_INIT_0F_BIT_00_C : bit_vector(255 downto 0) := x"4312DF2C54881EFCBD4494B9CA15F744750831230C3948536A0898E673695561";
   constant CPIX_NORMAL_INIT_0F_BIT_01_C : bit_vector(255 downto 0) := x"5BE0D4D01A1D49624F18D8ABEEAF67027831E7D9E8D1929941ED4C2463E150B8";
   constant CPIX_NORMAL_INIT_0F_BIT_02_C : bit_vector(255 downto 0) := x"94693564B3559281EB09563209AA3D8A0FA1AB0E0E2FB9FA857DCD838AFB8E81";
   constant CPIX_NORMAL_INIT_0F_BIT_03_C : bit_vector(255 downto 0) := x"FFE5C83D3E6847A29DCE5D50F101C382A99448DBEEC8D7402B594AB034AB7B06";
   constant CPIX_NORMAL_INIT_0F_BIT_04_C : bit_vector(255 downto 0) := x"0B47260C1F84034AEA9B0E4EEFA3D6293F0C17354358DB4E5E0513A52DC73ED6";
   constant CPIX_NORMAL_INIT_0F_BIT_05_C : bit_vector(255 downto 0) := x"1E352039042C5FA15B3961568A43D214900F1D2DBAC5A0972B38012723D363B4";
   constant CPIX_NORMAL_INIT_0F_BIT_06_C : bit_vector(255 downto 0) := x"2A7936152E914B78A4B121531675E7D6F4E7A96A9575730D20CC50150A7BC809";
   constant CPIX_NORMAL_INIT_0F_BIT_07_C : bit_vector(255 downto 0) := x"166B0DA4F80B45418F3BD5D2726F2A098C122F6282620FDF06397E78396BFDF3";
   constant CPIX_NORMAL_INIT_0F_BIT_08_C : bit_vector(255 downto 0) := x"546B1E4C66C05DF3754B33A9CE93F1EA5B9C41ED94334BA62F7465EE62C8874B";
   constant CPIX_NORMAL_INIT_0F_BIT_09_C : bit_vector(255 downto 0) := x"0CF30D787CD5AA9D7F55A72BE027A88061FD2C4A6D5FD0C2781B093C381A8AAB";
   constant CPIX_NORMAL_INIT_0F_BIT_10_C : bit_vector(255 downto 0) := x"0B75284D551991B7432D74C4CCF8AD57D09319043A7013FD4F6900AB0E220C2B";
   constant CPIX_NORMAL_INIT_0F_BIT_11_C : bit_vector(255 downto 0) := x"0919034C0E64AE73AE8C3A3C867E15F0C3411732B3F78454D0C37F2634665DF1";
   constant CPIX_NORMAL_INIT_0F_BIT_12_C : bit_vector(255 downto 0) := x"192A25255506C41E33925E3215F6B783B6122D203CEEBBB85D93FEAC3A3C0E04";
   constant CPIX_NORMAL_INIT_0F_BIT_13_C : bit_vector(255 downto 0) := x"056A425659981EF2C00653DB138C9D6F8D419793159CF1113F8FEE16A9995E23";
   constant CPIX_NORMAL_INIT_0F_BIT_14_C : bit_vector(255 downto 0) := x"103A8AE34341408969B1367F976789CF2B8DDB4E4BE5C7F346DEB26052CF42E9";
   constant CPIX_NORMAL_INIT_10_BIT_00_C : bit_vector(255 downto 0) := x"D30A96E9F18A9D98B10113A832B3033BB094764005BA8E9D50F2E0F4F752E986";
   constant CPIX_NORMAL_INIT_10_BIT_01_C : bit_vector(255 downto 0) := x"AB520B0CFF29C5B8D3807BC735492F66C29C4E1A6E5A67EA1350B7F5429CC5A1";
   constant CPIX_NORMAL_INIT_10_BIT_02_C : bit_vector(255 downto 0) := x"C31CF33ABDAD446686CE3942BEEB5723C878376C3FBBE9C5F6180B47C4B1167B";
   constant CPIX_NORMAL_INIT_10_BIT_03_C : bit_vector(255 downto 0) := x"722178AF942A1F961422BC3333D67360AF41E4A2DCD4AD35CE082E06A7FF1EC7";
   constant CPIX_NORMAL_INIT_10_BIT_04_C : bit_vector(255 downto 0) := x"BDFD399C877E7556B39CEE0246961CCBA4A96A9081E0266ED6CD73B6D759B0B6";
   constant CPIX_NORMAL_INIT_10_BIT_05_C : bit_vector(255 downto 0) := x"9B2BF0931829621BD33B35C53B6B31F3EAC447153B575C38C19B2206FB1995A9";
   constant CPIX_NORMAL_INIT_10_BIT_06_C : bit_vector(255 downto 0) := x"F31235231D99EE47C4015F3D2F80E64E03ED59287D0EC861CAEC5BFD845517C7";
   constant CPIX_NORMAL_INIT_10_BIT_07_C : bit_vector(255 downto 0) := x"8B7C16AF954D59CFE48A18D2D4FBBFFAF37FB61AED752D1D0B7A7CECAE863887";
   constant CPIX_NORMAL_INIT_10_BIT_08_C : bit_vector(255 downto 0) := x"669B76C1A21B93CE459508A1FA7F0BDBA93E049574E59C0F7E9A669F80FDAEFB";
   constant CPIX_NORMAL_INIT_10_BIT_09_C : bit_vector(255 downto 0) := x"1C012E5386D41F72ABBBB6405CD558220F24882511B34FB002ADF87C59B29EF5";
   constant CPIX_NORMAL_INIT_10_BIT_10_C : bit_vector(255 downto 0) := x"883A6D70C1A66EB319538D46745D32977233F9F7C20F130259FA0F34B3A8E7D4";
   constant CPIX_NORMAL_INIT_10_BIT_11_C : bit_vector(255 downto 0) := x"7EE463141B530B52C18541CDD55B2212B055B5EA40B1BA860B4B3351CBC7E87D";
   constant CPIX_NORMAL_INIT_10_BIT_12_C : bit_vector(255 downto 0) := x"0D97996C0C973A990D46C1B15A59C21585670326AFBE1DF514B464F0F2F81B51";
   constant CPIX_NORMAL_INIT_10_BIT_13_C : bit_vector(255 downto 0) := x"564DD8A5AF3A2DDC3EED386B19D39CEED7AB0541ED2CC79869FE435D5B60033D";
   constant CPIX_NORMAL_INIT_10_BIT_14_C : bit_vector(255 downto 0) := x"66FF1C6BF12BCEEBC5ADAF9716A398E98B19013C4A727B548725871E4D9ECB0C";
   constant CPIX_NORMAL_INIT_11_BIT_00_C : bit_vector(255 downto 0) := x"94495AD51C2EE5D441FDEB0CDAC85AEBC0FD3F4B22CB09ED592009BD4763C752";
   constant CPIX_NORMAL_INIT_11_BIT_01_C : bit_vector(255 downto 0) := x"D7D672294052F76DCE0866392DE7B229EAB8667174C89E3871113D8EDDD0EDFE";
   constant CPIX_NORMAL_INIT_11_BIT_02_C : bit_vector(255 downto 0) := x"79ED79B9F103CBD515DB91F136E337D21B6FB60194B2979CF4ABA2E4EC2B3492";
   constant CPIX_NORMAL_INIT_11_BIT_03_C : bit_vector(255 downto 0) := x"C9752AE352827D13324DB4E96631DFB00F62596E43787920ABC4CDD18780A71D";
   constant CPIX_NORMAL_INIT_11_BIT_04_C : bit_vector(255 downto 0) := x"49079E0245CC5C1B3EF214AFE7666B87329A7423133B34F25BDBCC4FCFAB0A4E";
   constant CPIX_NORMAL_INIT_11_BIT_05_C : bit_vector(255 downto 0) := x"93D6A14541D76F168B98BA3E08906A1635734C4869D0277AC6F5D2F0191D9AE6";
   constant CPIX_NORMAL_INIT_11_BIT_06_C : bit_vector(255 downto 0) := x"74598E34976A98B6356D8582539D880FFDF1E6155AFB3135A19B672C6267978D";
   constant CPIX_NORMAL_INIT_11_BIT_07_C : bit_vector(255 downto 0) := x"8878417B5E42A8099F4F2626D74B78ED81C806E963EA04B3571A58C22E6AC1CA";
   constant CPIX_NORMAL_INIT_11_BIT_08_C : bit_vector(255 downto 0) := x"A3A6CC407DA5F3983F808F3537E6B882A4BC63131D634B460E4BEC1B9E5BF30D";
   constant CPIX_NORMAL_INIT_11_BIT_09_C : bit_vector(255 downto 0) := x"5DC046DC7058CB1D42548F71EF2B6D438269679966677F9D3DE3B7965EF67C99";
   constant CPIX_NORMAL_INIT_11_BIT_10_C : bit_vector(255 downto 0) := x"4F25EF003E2247D5777A666C036982D64B231F2552F717F3904BB775FFF611B7";
   constant CPIX_NORMAL_INIT_11_BIT_11_C : bit_vector(255 downto 0) := x"41373DAB70015CF428ABF77FF355ED787F55424AA722B2A725ACC81D06F2F11E";
   constant CPIX_NORMAL_INIT_11_BIT_12_C : bit_vector(255 downto 0) := x"89FECBEC45BC2358A3A3D0FA6BC4C37DE457F681DDE7438BB1FD00D35B531363";
   constant CPIX_NORMAL_INIT_11_BIT_13_C : bit_vector(255 downto 0) := x"1F3A3F969D46C21FA7533A5A121C1C47692BDE4038B8A8FCDD80C9B0DE42A897";
   constant CPIX_NORMAL_INIT_11_BIT_14_C : bit_vector(255 downto 0) := x"C07821686940C2B233344BCCFB7DA96512BAA9670004E96FD1B503D11E8796BD";
   constant CPIX_NORMAL_INIT_12_BIT_00_C : bit_vector(255 downto 0) := x"0DF38DECC4DE0C4C3B32D0B94155C3015A2AF491BB0B469146B59F6E54521A23";
   constant CPIX_NORMAL_INIT_12_BIT_01_C : bit_vector(255 downto 0) := x"F5E86592D3FB8390B2CAB679CD6FC268C25DE819D944E09C5F583B7CE205B128";
   constant CPIX_NORMAL_INIT_12_BIT_02_C : bit_vector(255 downto 0) := x"E5F50B5F8816130D9BE79F6329CF6AD0FC60684DADEE66ABE60610FD8E7DD7EC";
   constant CPIX_NORMAL_INIT_12_BIT_03_C : bit_vector(255 downto 0) := x"FCD1930D6E72D1EA427B7F2207C903A595CA44CC4F2EE6AB0DA3366D2DEB9E2E";
   constant CPIX_NORMAL_INIT_12_BIT_04_C : bit_vector(255 downto 0) := x"1C651BD421D9A47EFFD72E008DFD8480D6C38DF0BCCAFCA027E0FFACF3878297";
   constant CPIX_NORMAL_INIT_12_BIT_05_C : bit_vector(255 downto 0) := x"60990BE498FC7EF1594AF92452A080154E5A091947A337FAC175D552B9EA9D4E";
   constant CPIX_NORMAL_INIT_12_BIT_06_C : bit_vector(255 downto 0) := x"923AFF8B52B4B1CF38C117F88702DE415123464DEEB0A005DB8CCF42EC30A836";
   constant CPIX_NORMAL_INIT_12_BIT_07_C : bit_vector(255 downto 0) := x"1C0BC6AFD95AE648EB3E25A8895FED28468B72408C440086588A01E06A3F7562";
   constant CPIX_NORMAL_INIT_12_BIT_08_C : bit_vector(255 downto 0) := x"6AD763F306FF68927E2F3EB3F45D9986FC9CB11755BEFF730B9A581E664D5AD5";
   constant CPIX_NORMAL_INIT_12_BIT_09_C : bit_vector(255 downto 0) := x"CAF9CCD8438B87DC6CD5DFB45B8FBB17DA74E5FE517BDFF99D5013BF976E0D3F";
   constant CPIX_NORMAL_INIT_12_BIT_10_C : bit_vector(255 downto 0) := x"E2F3482B0F7BBF6495444A795A3F66D0D46EBA9B469DB71B09C12FBF51CFF2D9";
   constant CPIX_NORMAL_INIT_12_BIT_11_C : bit_vector(255 downto 0) := x"F7B5FAF464FA458F3B24EC5CEC1F58FBB9EABDB1F497BF596B3DC2179D0DE631";
   constant CPIX_NORMAL_INIT_12_BIT_12_C : bit_vector(255 downto 0) := x"7852EC947C4DE48E60729D9364BD356692AFBB58D876BF55453168DE671D07DF";
   constant CPIX_NORMAL_INIT_12_BIT_13_C : bit_vector(255 downto 0) := x"53BB3F1EC03B1884CED2C4F82D2D5AAFD324659AF6529FD1F97E2D99A5AE8159";
   constant CPIX_NORMAL_INIT_12_BIT_14_C : bit_vector(255 downto 0) := x"9898FCE1FC372C6150F8F076E607CE0E1F07A2B9ECF0971741CCC0DB681A5714";
   constant CPIX_NORMAL_INIT_13_BIT_00_C : bit_vector(255 downto 0) := x"D50CBEE6ACFA27DA9B52891B65B607D0A50B8D2F7BA9509485D51D4470795465";
   constant CPIX_NORMAL_INIT_13_BIT_01_C : bit_vector(255 downto 0) := x"E070B6C74614DB3455864D0898A70EC9B950944140E8BF93005D1DF48C3ED7DE";
   constant CPIX_NORMAL_INIT_13_BIT_02_C : bit_vector(255 downto 0) := x"60637D0C6DD875876AA9ACF73B7F1FDED1E4269565B38641F155C7DD00BBC0AC";
   constant CPIX_NORMAL_INIT_13_BIT_03_C : bit_vector(255 downto 0) := x"8C5D2A6C54F0EF519664B3C53742DF0D2C89F341573CC8CC5B73A766267DC61D";
   constant CPIX_NORMAL_INIT_13_BIT_04_C : bit_vector(255 downto 0) := x"82D28BE4277EBA4B9289404963EC97D7D5F20B4C5DFF2A72BE92155B3A032B0A";
   constant CPIX_NORMAL_INIT_13_BIT_05_C : bit_vector(255 downto 0) := x"F3D4EF331C925D49818AAEFA72E919CE4DCE878F9B8166D10DC163BDBC8C4E52";
   constant CPIX_NORMAL_INIT_13_BIT_06_C : bit_vector(255 downto 0) := x"8A3680F62A27C9D00DBAD9E9EDA0FA9EED380C44C9F9FB67AE30A5023E98867A";
   constant CPIX_NORMAL_INIT_13_BIT_07_C : bit_vector(255 downto 0) := x"A819A324E95D9B8BD580AE68564F927583B3D9F28C6EFA41439AE925E7A1A9A1";
   constant CPIX_NORMAL_INIT_13_BIT_08_C : bit_vector(255 downto 0) := x"DD19D1B131D88DE83BC96F19935F2DC834085E7C64E664BB8FCF08D187B31B7E";
   constant CPIX_NORMAL_INIT_13_BIT_09_C : bit_vector(255 downto 0) := x"BCF5881DB2C93A6DCAD47E934C592F44F679B345C23A81939C5178371AB2D68C";
   constant CPIX_NORMAL_INIT_13_BIT_10_C : bit_vector(255 downto 0) := x"3372613B49DF260A857BD026BDDBFD4A3823B350502C7160DEE1C8BE3AC6FE59";
   constant CPIX_NORMAL_INIT_13_BIT_11_C : bit_vector(255 downto 0) := x"91AC38B75B0E4D9B50723B6B51EBBEAA3FA73DDA537988D61F8732B8ED28E5B0";
   constant CPIX_NORMAL_INIT_13_BIT_12_C : bit_vector(255 downto 0) := x"9745C1302E6AFEA7BD46950998DBB2BA330A1A33BBA0BA5CE6FB6BB19DE4CAE8";
   constant CPIX_NORMAL_INIT_13_BIT_13_C : bit_vector(255 downto 0) := x"9AF027FB68E31BB04E8572A765F94E85673F9064ADD5A95C90C6E013BC2C19C3";
   constant CPIX_NORMAL_INIT_13_BIT_14_C : bit_vector(255 downto 0) := x"22A52A5BBD725E1789A5E0ECAD5ABA9B174259A4A26F77639D4EFFF251C3EA16";
   constant CPIX_NORMAL_INIT_14_BIT_00_C : bit_vector(255 downto 0) := x"7C2779BFD4D894211FC73045F06952CFEA0172B29FFAE1203BFD9F58595A56CE";
   constant CPIX_NORMAL_INIT_14_BIT_01_C : bit_vector(255 downto 0) := x"6E77D97C08883F33B29AAFC1E230409FB518785052FF77E9B3EA69B8C9F879ED";
   constant CPIX_NORMAL_INIT_14_BIT_02_C : bit_vector(255 downto 0) := x"D9727B86A337C986538F58D8A86E4425B08ABBE0DE69C41B39855933560EEE56";
   constant CPIX_NORMAL_INIT_14_BIT_03_C : bit_vector(255 downto 0) := x"2E6CC3CFF3DA7881B308ABC263DDF426235149AB4F60E3549BF1BF8BC1D904F7";
   constant CPIX_NORMAL_INIT_14_BIT_04_C : bit_vector(255 downto 0) := x"3C07C56C1BD72C685D06F61C45B5C3AD9347C621CFD1F3A5D0C405220A262CA2";
   constant CPIX_NORMAL_INIT_14_BIT_05_C : bit_vector(255 downto 0) := x"E8FBA852ABEB3E14743053C156820BD3BDA0E687AFAA0249C72AEC9527D92DDD";
   constant CPIX_NORMAL_INIT_14_BIT_06_C : bit_vector(255 downto 0) := x"FCC588CAEED47B3E614821880428BF69FD9DAC9C53989B48E1704B20E848A37F";
   constant CPIX_NORMAL_INIT_14_BIT_07_C : bit_vector(255 downto 0) := x"D14BED2114AEC096A5116BB5D999305CF3101C00DFB12ADEE08A19AB77E36B87";
   constant CPIX_NORMAL_INIT_14_BIT_08_C : bit_vector(255 downto 0) := x"187D1A3DC17280CA02D9A5B5B3F147F5B4C46F3495C10D319DE462CB269FDDA6";
   constant CPIX_NORMAL_INIT_14_BIT_09_C : bit_vector(255 downto 0) := x"EDF60731BA6C1B1FFAA5AB22DAF41EB6FE8254FBFC065318E303CFBC84F0BA96";
   constant CPIX_NORMAL_INIT_14_BIT_10_C : bit_vector(255 downto 0) := x"A8B581DADCAA92A5810213937AD79E3CEA321B8F2FBEDB0699BB489043670E2F";
   constant CPIX_NORMAL_INIT_14_BIT_11_C : bit_vector(255 downto 0) := x"BA5CF46FDE1BC6CC65406D581E97F87F8EBB4952DA0AE1E2B112FEB033ECB334";
   constant CPIX_NORMAL_INIT_14_BIT_12_C : bit_vector(255 downto 0) := x"047F778C65F02CC3DC0C309E925B2FD802E795FB44572552CED7746EEA98FE4E";
   constant CPIX_NORMAL_INIT_14_BIT_13_C : bit_vector(255 downto 0) := x"8F877C85BFD9A89C82AF1DEF7CD028B80BDFA73A5E87DAC47E4FFA4F18BD5532";
   constant CPIX_NORMAL_INIT_14_BIT_14_C : bit_vector(255 downto 0) := x"B638D6270696952B4A07EC27A55813FA7DB48F8E133F952DEE6F27069779B706";
   constant CPIX_NORMAL_INIT_15_BIT_00_C : bit_vector(255 downto 0) := x"7899A1E62739A82395BC81225AF08975EA095287B11DD152CA3305EA86D353ED";
   constant CPIX_NORMAL_INIT_15_BIT_01_C : bit_vector(255 downto 0) := x"44F3F7F16B1A9F0B4C082A6D2C7114D59E692A9CD0470531CB85555D1451B873";
   constant CPIX_NORMAL_INIT_15_BIT_02_C : bit_vector(255 downto 0) := x"49CDF24D63EA682A8AE08932F6784A54CD34D30EB00F2DB3FBE1CFF9F50BFE0B";
   constant CPIX_NORMAL_INIT_15_BIT_03_C : bit_vector(255 downto 0) := x"937B8E7A51832F959844EE153343839717D0DFCC350C09D4671BA566C20F5CB7";
   constant CPIX_NORMAL_INIT_15_BIT_04_C : bit_vector(255 downto 0) := x"301BD97EF1B9E219DD00D811EAF9C3D4AD23119A30CDA1A6C22DDCEEEF440FC6";
   constant CPIX_NORMAL_INIT_15_BIT_05_C : bit_vector(255 downto 0) := x"C9D007B39B85193B6663C40B744F6E28F6DC973237BA35D18D877984055F6CA7";
   constant CPIX_NORMAL_INIT_15_BIT_06_C : bit_vector(255 downto 0) := x"A0669B3F784ACA4F360BEC814ACAD81AE20EA71CCABE747EF6DA987376EFC309";
   constant CPIX_NORMAL_INIT_15_BIT_07_C : bit_vector(255 downto 0) := x"15365A0EF225DDD849D1B4D51B3A72CFAF0B7EEBCEF4CAB23B8310CFFFA56140";
   constant CPIX_NORMAL_INIT_15_BIT_08_C : bit_vector(255 downto 0) := x"6DD139F698527EE04A875F8FF5B45614E8285EF55753D1A3F904F55182C3DBF6";
   constant CPIX_NORMAL_INIT_15_BIT_09_C : bit_vector(255 downto 0) := x"E0FBFA88DFB08C2B945B2E70A7BC40BCF4D18BF15B9A31D995293EDC8F9703C6";
   constant CPIX_NORMAL_INIT_15_BIT_10_C : bit_vector(255 downto 0) := x"D9EE231A6156EE5B28344D648E13E9A9EB780E47728CF3A5ACD5FE1ED34BC2D0";
   constant CPIX_NORMAL_INIT_15_BIT_11_C : bit_vector(255 downto 0) := x"E320D0B4FBCD709BED8793696BF0028EBCB175ED979140CB29F26CB496FD6D0C";
   constant CPIX_NORMAL_INIT_15_BIT_12_C : bit_vector(255 downto 0) := x"82FE7B8CE5E80F666E91DA5BA1A7530DD30666913652E97C3906C2970B4CBE5C";
   constant CPIX_NORMAL_INIT_15_BIT_13_C : bit_vector(255 downto 0) := x"34B0456B9ED21A4CFE7C6851A1EF94C7FE796884C7136B803E3430187DE7C022";
   constant CPIX_NORMAL_INIT_15_BIT_14_C : bit_vector(255 downto 0) := x"041B0C38C90724E29119F0B07D86CDA27839B9D3244B85892C9E57F6E57CBDED";
   constant CPIX_NORMAL_INIT_16_BIT_00_C : bit_vector(255 downto 0) := x"C12AFD7BBE881FBD8F0F92A7EEADEABF50D99E7A44ACB9D19E4A94FB6EE27BF0";
   constant CPIX_NORMAL_INIT_16_BIT_01_C : bit_vector(255 downto 0) := x"507ADB6BB621EDE35CB2A3525E81D0C625519211CF876EE2E1441C8B25093A7D";
   constant CPIX_NORMAL_INIT_16_BIT_02_C : bit_vector(255 downto 0) := x"8CF54BB1383175F73AFF14C81C4BAF5C1FC62EF6B3D06A0EBE13CF16E6ECE0D1";
   constant CPIX_NORMAL_INIT_16_BIT_03_C : bit_vector(255 downto 0) := x"3AFB3A297FFA7441AEFC172D6710234A7898E791ABAFB5C77B93DFCA4A75BE04";
   constant CPIX_NORMAL_INIT_16_BIT_04_C : bit_vector(255 downto 0) := x"804E3AACA724295C78B2C2C514AA10FB156FD849861B8D9F849DD8BF6AF697E1";
   constant CPIX_NORMAL_INIT_16_BIT_05_C : bit_vector(255 downto 0) := x"30E20EB9F8E24E6D36599324D8992CA22098969C1510384176BC70BFDD0EACDF";
   constant CPIX_NORMAL_INIT_16_BIT_06_C : bit_vector(255 downto 0) := x"63F08F9BEB85BD42DC80B6E78B5085C2F441717185A2A2B5999046C7D9BA9252";
   constant CPIX_NORMAL_INIT_16_BIT_07_C : bit_vector(255 downto 0) := x"B41861DEF4E0E4142474EF8B37C579C45358DB2D8BD498498A1E04867847464F";
   constant CPIX_NORMAL_INIT_16_BIT_08_C : bit_vector(255 downto 0) := x"204947682E95F04DD5D05C82965DBF13A8959562B0EE2343B9048D52AFCF76E7";
   constant CPIX_NORMAL_INIT_16_BIT_09_C : bit_vector(255 downto 0) := x"891D23430264BD53152B22731B4E3F90D7A80540E011B7931F5E489135DFAF4D";
   constant CPIX_NORMAL_INIT_16_BIT_10_C : bit_vector(255 downto 0) := x"ECC6292A5D5C3B776E947B5F77E8F7DB5C6291B7D7725177EC9DB666E1388B22";
   constant CPIX_NORMAL_INIT_16_BIT_11_C : bit_vector(255 downto 0) := x"257E7A0FE83784CB9550591C9F42F9AEAD90EB0A4DB88D5CD660010C925E555C";
   constant CPIX_NORMAL_INIT_16_BIT_12_C : bit_vector(255 downto 0) := x"2F70F2955A9ECE88681023E6D676E11256D5D9E96C9D098A914C0C817490320B";
   constant CPIX_NORMAL_INIT_16_BIT_13_C : bit_vector(255 downto 0) := x"329D468301CA664F2B6FD393DA40D55FA1CB865B712D68899C074084AD1FC488";
   constant CPIX_NORMAL_INIT_16_BIT_14_C : bit_vector(255 downto 0) := x"96DA7CF176D425E8E66E10516C729BBA6CE8FACE931F646769F3FB6E436FEBB8";
   constant CPIX_NORMAL_INIT_17_BIT_00_C : bit_vector(255 downto 0) := x"D333BB1B89CD1C43AC85410C5CD6CD6FE7FC7B10060E1E2D62CE6B530440FF9D";
   constant CPIX_NORMAL_INIT_17_BIT_01_C : bit_vector(255 downto 0) := x"CBC5A282E29C95D597BB5508E65485A14A07A05FCF337FF0BF2865A5680384BA";
   constant CPIX_NORMAL_INIT_17_BIT_02_C : bit_vector(255 downto 0) := x"0B0D4394760C2966E96F2A0A9535384976BB708A0175120D11C53043E1C6E539";
   constant CPIX_NORMAL_INIT_17_BIT_03_C : bit_vector(255 downto 0) := x"E4CBC0DB50E78B9061611B0524E42D4E18868DB1DDA4FCCF031A0A17882EF3F4";
   constant CPIX_NORMAL_INIT_17_BIT_04_C : bit_vector(255 downto 0) := x"9DBC38DB5AC1268C17CABCD9A9D6AB85EB0542153F4B9B07DF9B28F050ACC041";
   constant CPIX_NORMAL_INIT_17_BIT_05_C : bit_vector(255 downto 0) := x"A97E392E0E3D02E9DCB1C71B17E6A38964A4A2E25FA71F8F189CBDE420CFE366";
   constant CPIX_NORMAL_INIT_17_BIT_06_C : bit_vector(255 downto 0) := x"9EEA025C2F8D77C74EA557FA1469DE7EB2747ED1F3DA92083C04A5E3BB151AFC";
   constant CPIX_NORMAL_INIT_17_BIT_07_C : bit_vector(255 downto 0) := x"8AEDA4DE11DC0CC2A9ABA48AB82617B256D46FE8E81994B0F7069962D473B5D1";
   constant CPIX_NORMAL_INIT_17_BIT_08_C : bit_vector(255 downto 0) := x"03F299477A481061D13642F1ADB0D8B6AB7671AD6A68921B9255BA96A84AD958";
   constant CPIX_NORMAL_INIT_17_BIT_09_C : bit_vector(255 downto 0) := x"1A1FA04F9001F90C78F9903E9A2328FE51D90B663654A42EDEDD24B278CEEFC0";
   constant CPIX_NORMAL_INIT_17_BIT_10_C : bit_vector(255 downto 0) := x"7C779EA4C4021D65BED0349DEB6C3330A4FA202AB6040D4D2D20F86C5FEDFBF2";
   constant CPIX_NORMAL_INIT_17_BIT_11_C : bit_vector(255 downto 0) := x"581A3B3283DB7A5C5E835E9F8A5602D63DF4725039E15A499570F75AC55B220A";
   constant CPIX_NORMAL_INIT_17_BIT_12_C : bit_vector(255 downto 0) := x"46B37791D321214389B4A63EC5E3588C551FDAA559DF8F4F9486CF592F5C8FCD";
   constant CPIX_NORMAL_INIT_17_BIT_13_C : bit_vector(255 downto 0) := x"48116FD06284755E7E6E59DE384C16BFA88878F41298B4FE2FAFE956961057C7";
   constant CPIX_NORMAL_INIT_17_BIT_14_C : bit_vector(255 downto 0) := x"1C8C6C34B98DEEE4B44629B992A4646C5793B458BBBA4E65D637F8674F8A093C";
   constant CPIX_NORMAL_INIT_18_BIT_00_C : bit_vector(255 downto 0) := x"7DA1CB0438FF571E776A8D69AA5594E9FAC75B6FBA09F9F09ECD4C18776EDBA1";
   constant CPIX_NORMAL_INIT_18_BIT_01_C : bit_vector(255 downto 0) := x"4B446566AB427E16518A15FE3F858CA961F6105FF690ACE1A3972083C054C76B";
   constant CPIX_NORMAL_INIT_18_BIT_02_C : bit_vector(255 downto 0) := x"3A52FED6D47105A6921480436857E40B00E5481B42309D9B6E308BB3052E767C";
   constant CPIX_NORMAL_INIT_18_BIT_03_C : bit_vector(255 downto 0) := x"866036C3AF1AB50EA6FB05ED0D30784AA1AE064F8F57394611431532A3C4A57D";
   constant CPIX_NORMAL_INIT_18_BIT_04_C : bit_vector(255 downto 0) := x"658BBB5D3B0F3F2703635F78548255C6305718C05DC096DC41868A4B2B35F723";
   constant CPIX_NORMAL_INIT_18_BIT_05_C : bit_vector(255 downto 0) := x"B040363DFBF4C94FFEC0218610574AF2C27A68239C19DE2021946FFE7FEAD5A6";
   constant CPIX_NORMAL_INIT_18_BIT_06_C : bit_vector(255 downto 0) := x"6BA0B9DB1D9C5187BA858412FECD2D08BD8381682CDB79872793F774B66AFB87";
   constant CPIX_NORMAL_INIT_18_BIT_07_C : bit_vector(255 downto 0) := x"DCDD92AC2378D779B360D5450D21859EB72A56A032AF6015B765B7040DE86F9C";
   constant CPIX_NORMAL_INIT_18_BIT_08_C : bit_vector(255 downto 0) := x"FA2DA1210BD9F694BE0418D20564DC1D860B853495EA75D4841331F9961211E6";
   constant CPIX_NORMAL_INIT_18_BIT_09_C : bit_vector(255 downto 0) := x"EC60EF1A124C19AC3268D2F18D8D1F2F98F56E7B21F5DC4BB9850CA39797834F";
   constant CPIX_NORMAL_INIT_18_BIT_10_C : bit_vector(255 downto 0) := x"270B3C529582B80C991DA8CFAED8FDCBB734FBBE9C731FAFADD207961F094955";
   constant CPIX_NORMAL_INIT_18_BIT_11_C : bit_vector(255 downto 0) := x"3B57FFED9B1F85190EC69B09BDEAA78455B1FAAFCE17EE9052C4DC316D2604A5";
   constant CPIX_NORMAL_INIT_18_BIT_12_C : bit_vector(255 downto 0) := x"77ED6A1F543325DBF090D0C8473EE60F95FA6A8B33C03F8873B97A4F7DAF630F";
   constant CPIX_NORMAL_INIT_18_BIT_13_C : bit_vector(255 downto 0) := x"91EDF87EFCFA86EC2224BB21D9DB8C6F80ED6F1FF06D09FC1856EBC4E3445656";
   constant CPIX_NORMAL_INIT_18_BIT_14_C : bit_vector(255 downto 0) := x"06184CB647EE647F163B098FE464BAF6B4791B2EDBA6B86CA0EBE210603D1A6A";
   constant CPIX_NORMAL_INIT_19_BIT_00_C : bit_vector(255 downto 0) := x"CEB4975BF10BFE85076B9C85DF009D0E1BB37A6E2806B825F3CDF05EB0435072";
   constant CPIX_NORMAL_INIT_19_BIT_01_C : bit_vector(255 downto 0) := x"64D5DDB7770CB94B637372D5E19E57311F3D3AB6DB9694906D57C6089E773375";
   constant CPIX_NORMAL_INIT_19_BIT_02_C : bit_vector(255 downto 0) := x"07347EB0A01640077FAD604B344C8EE4DD7E6831FD68FECC8A8B7B44F484C494";
   constant CPIX_NORMAL_INIT_19_BIT_03_C : bit_vector(255 downto 0) := x"987B2299F8AC3E296063158F209870815E0E5664A9857FE9312CDDBBE303F86B";
   constant CPIX_NORMAL_INIT_19_BIT_04_C : bit_vector(255 downto 0) := x"12045A9FD95D50B7307F600C210F97B1C0266299A187A0AD21A4C6FC9E56779A";
   constant CPIX_NORMAL_INIT_19_BIT_05_C : bit_vector(255 downto 0) := x"E164444EFA7A21BEFB5B4E3966A148B76EB2196BEEFB3A6774DB50B590D84451";
   constant CPIX_NORMAL_INIT_19_BIT_06_C : bit_vector(255 downto 0) := x"F5CAD74A7C795BC1854F5D5CCFE7272EFF4E5DA4AC5A83C00ACF07666CC53F23";
   constant CPIX_NORMAL_INIT_19_BIT_07_C : bit_vector(255 downto 0) := x"87F76F204D2957BE98C68779F7EE97CF15D9BE0534E268620E22D5A12E5A6B76";
   constant CPIX_NORMAL_INIT_19_BIT_08_C : bit_vector(255 downto 0) := x"B1ED24E073763F10F0308745567E1BFA02006F47B76405FB95FA2EB26EAEC87D";
   constant CPIX_NORMAL_INIT_19_BIT_09_C : bit_vector(255 downto 0) := x"13C646539F5449E50750EE576E2FC356003D19DB1E8EC1E687895C5BC77FF691";
   constant CPIX_NORMAL_INIT_19_BIT_10_C : bit_vector(255 downto 0) := x"353568F6341A11AAD57EB4E1AEA3E3BEFCBAABAC164C21211B0939B4FC565605";
   constant CPIX_NORMAL_INIT_19_BIT_11_C : bit_vector(255 downto 0) := x"0FE18AB9D7577A92BC4005ABAE965BB70C8E9AB908E77E8411CBB67355AA8240";
   constant CPIX_NORMAL_INIT_19_BIT_12_C : bit_vector(255 downto 0) := x"1C923B0622D29DA2B779747E9E8CB392C69F92A63861F97DBC0A771B20E0A8BC";
   constant CPIX_NORMAL_INIT_19_BIT_13_C : bit_vector(255 downto 0) := x"3DA560304406A24879DBA4EDA6143141591B514BE9AAE6694BA24E76E94AB9F0";
   constant CPIX_NORMAL_INIT_19_BIT_14_C : bit_vector(255 downto 0) := x"1BCB42567EFA469B82B044453611FA80D9DAFA90D33FF6DF329C73B10003DE0E";
   constant CPIX_NORMAL_INIT_1A_BIT_00_C : bit_vector(255 downto 0) := x"7E40EB0403DA24E64F1BC4F48B5CFB2315C2788EF8D97974AA51BE40D18FDCF2";
   constant CPIX_NORMAL_INIT_1A_BIT_01_C : bit_vector(255 downto 0) := x"F1FE2E454E9724AE18AC5A777E37D92EED604D73A362A6E2DBD81C9631AEA60F";
   constant CPIX_NORMAL_INIT_1A_BIT_02_C : bit_vector(255 downto 0) := x"CCA0E37A127F5DA12E14AEB3FF0E5D87AC3A999DD5E6C5D29A1E4F5462D011A0";
   constant CPIX_NORMAL_INIT_1A_BIT_03_C : bit_vector(255 downto 0) := x"89085C9CCFF1D5419965EE191014AE9F24740CAA90D99BC2935C45ECF0BDE1B1";
   constant CPIX_NORMAL_INIT_1A_BIT_04_C : bit_vector(255 downto 0) := x"83400DB7DC59090DB81203DE58FED07BF12373A6906938CBAB1A1712C72714E6";
   constant CPIX_NORMAL_INIT_1A_BIT_05_C : bit_vector(255 downto 0) := x"BBB6CC18B26319AE5F67D4C7CEA5C9974215D08744F4BF44F2346299EA8F4E73";
   constant CPIX_NORMAL_INIT_1A_BIT_06_C : bit_vector(255 downto 0) := x"9AFC84EAD905C68A3DD8F712B86D465A923414795AE55D1FE9555C8DCA983013";
   constant CPIX_NORMAL_INIT_1A_BIT_07_C : bit_vector(255 downto 0) := x"3DC6412793FCE09261B19F83D77435827831DCD53E4DB5806015026C2ACC2D95";
   constant CPIX_NORMAL_INIT_1A_BIT_08_C : bit_vector(255 downto 0) := x"EE355043C075018C9217DFA70EBBDFCC8074546BAB96CA6075091E765828F6F5";
   constant CPIX_NORMAL_INIT_1A_BIT_09_C : bit_vector(255 downto 0) := x"B79A2DC80D2DF903EF05FF5F774A9ACFB169CF282A2D2770D8040575648097D7";
   constant CPIX_NORMAL_INIT_1A_BIT_10_C : bit_vector(255 downto 0) := x"44BD4BBBEE02ECCA88CBD7205BD4212485D53F330ECEA1BF227B9BAF09C625AD";
   constant CPIX_NORMAL_INIT_1A_BIT_11_C : bit_vector(255 downto 0) := x"6B548B16630E53F741D696981BAB2732B4272B4C976662CFBEFFA3B64FFF9727";
   constant CPIX_NORMAL_INIT_1A_BIT_12_C : bit_vector(255 downto 0) := x"FA493F155D83DE1639A7954A682D6901FA46FF90968AD68EA6FA6597D7BA21AA";
   constant CPIX_NORMAL_INIT_1A_BIT_13_C : bit_vector(255 downto 0) := x"DD2519209E73AB53927A2DB66B79A8325CAF9F27D4868B9367FE2DBA1297ED68";
   constant CPIX_NORMAL_INIT_1A_BIT_14_C : bit_vector(255 downto 0) := x"B9231F46C8E6996EEBBE554293D1B3FF0A7C5F16413330F72A7F5FE3298AB4FC";
   constant CPIX_NORMAL_INIT_1B_BIT_00_C : bit_vector(255 downto 0) := x"C8F0C23DD066192359957DD30D104FE4AA9B57F3E72C7A8116392BD7E565862F";
   constant CPIX_NORMAL_INIT_1B_BIT_01_C : bit_vector(255 downto 0) := x"53331F8B4D85513892463A652F75258499DBBDA5451FB4AB9B2A41B88D268D5A";
   constant CPIX_NORMAL_INIT_1B_BIT_02_C : bit_vector(255 downto 0) := x"079C1AC0F351616F134E5035135F1178B007FD72D341555459FC5232FC2E90C9";
   constant CPIX_NORMAL_INIT_1B_BIT_03_C : bit_vector(255 downto 0) := x"F90071D2F2BBA575559AEF6DB6E547F6BE9834132914BA75A5B2AFAEC6B8C0A9";
   constant CPIX_NORMAL_INIT_1B_BIT_04_C : bit_vector(255 downto 0) := x"50F7A41BEAD0E5F6B251F3750B2DF0AE6285C5645AE6B692EEFC0D645FBA8A17";
   constant CPIX_NORMAL_INIT_1B_BIT_05_C : bit_vector(255 downto 0) := x"67F9856258B4E77B1715A969BE3C9749124B8EE3845C1F181E62C10D9CF6B879";
   constant CPIX_NORMAL_INIT_1B_BIT_06_C : bit_vector(255 downto 0) := x"1595780F3ED183B3A923165F18E8A7ED280D4666DB3BE1894F12A7A5647DC205";
   constant CPIX_NORMAL_INIT_1B_BIT_07_C : bit_vector(255 downto 0) := x"564A81CCA944371FBE609BBCC309D21634F606D9F08DC096B3F19FD70E2E96A8";
   constant CPIX_NORMAL_INIT_1B_BIT_08_C : bit_vector(255 downto 0) := x"444DBC144F15E68EA28E230B73806249EBF46033755475C889FC317D10B741C6";
   constant CPIX_NORMAL_INIT_1B_BIT_09_C : bit_vector(255 downto 0) := x"111B93D92994F1C2E0D35D72BF636D3B50473E396108777409BF6202E9D68111";
   constant CPIX_NORMAL_INIT_1B_BIT_10_C : bit_vector(255 downto 0) := x"A5E99EFDF289A62DA086BEE94B67F655D9037FD907A3FF9786146DD72E2E2865";
   constant CPIX_NORMAL_INIT_1B_BIT_11_C : bit_vector(255 downto 0) := x"2563F89417971C15D6C0DC6FA83F517DEAABFD953BD380739BBF2890DA2A9A4A";
   constant CPIX_NORMAL_INIT_1B_BIT_12_C : bit_vector(255 downto 0) := x"6E827176AEE7F55C2145ED05576236C282482D70962F7DAA2DC0713FC2C3FE9F";
   constant CPIX_NORMAL_INIT_1B_BIT_13_C : bit_vector(255 downto 0) := x"22795567A67294D685AF7A51BAB7DFF37D69AE1369EB868E4C199149471D0703";
   constant CPIX_NORMAL_INIT_1B_BIT_14_C : bit_vector(255 downto 0) := x"45C8E03E8BF83BB5805C014CAE4EB32C4D96E01457A367BA1927BB6460BC8948";
   constant CPIX_NORMAL_INIT_1C_BIT_00_C : bit_vector(255 downto 0) := x"9F6606553E21DC84A4F4EE889C2E42FCDE745B30B88E826328E85E27B8B23DBA";
   constant CPIX_NORMAL_INIT_1C_BIT_01_C : bit_vector(255 downto 0) := x"8F892B6C06AF7F4D347E730F12D0976A595297964B18700AD6B1FBCBA5DD174E";
   constant CPIX_NORMAL_INIT_1C_BIT_02_C : bit_vector(255 downto 0) := x"D51E88A68F9BBF23FC366F63354245AF64684491C66D6D4B870221A3227F70D0";
   constant CPIX_NORMAL_INIT_1C_BIT_03_C : bit_vector(255 downto 0) := x"A30E2DAE9FD55F800C97D7B4C6BBE9F29AD0231FC5288884D5948EDE46BF61F9";
   constant CPIX_NORMAL_INIT_1C_BIT_04_C : bit_vector(255 downto 0) := x"60BB84FD69453E2C789F526ED8FC33259DE0C17F1D2C0D2F527B4D9E9670D194";
   constant CPIX_NORMAL_INIT_1C_BIT_05_C : bit_vector(255 downto 0) := x"A9DEA85C8665F9F999F6FBE19A6BCF3C0DED4018B433DCCD949FE76977BA3FE0";
   constant CPIX_NORMAL_INIT_1C_BIT_06_C : bit_vector(255 downto 0) := x"12F7468B51B7E715948E91C30420EC2B97F1941932461038F8EFAADFB3FCD468";
   constant CPIX_NORMAL_INIT_1C_BIT_07_C : bit_vector(255 downto 0) := x"6B787CFCEAD4BDE3C97B24815454FDFE956C00B1EC6CD643279855F1A4994271";
   constant CPIX_NORMAL_INIT_1C_BIT_08_C : bit_vector(255 downto 0) := x"BA4E4AD18E48D654CFB7C5FE76D11735E303F0A930974E395292E80C186B4042";
   constant CPIX_NORMAL_INIT_1C_BIT_09_C : bit_vector(255 downto 0) := x"4A92072C3918E1EC2F51A8D1FAAFEF70ECE63C4A9CD4723D63BC0F00E89D460D";
   constant CPIX_NORMAL_INIT_1C_BIT_10_C : bit_vector(255 downto 0) := x"79055239903F2516B9DCCB11F3EB3712965372FE7D90A3DAC53123A87CC01243";
   constant CPIX_NORMAL_INIT_1C_BIT_11_C : bit_vector(255 downto 0) := x"C0B28612A4A7E6B25FB353A1344819DB5F23B31ABA3DFECB51477B829DA3F02E";
   constant CPIX_NORMAL_INIT_1C_BIT_12_C : bit_vector(255 downto 0) := x"7505A8107B8A658C159AC5DEF3E49F3914ABFBDBCCAD1B21B3A470F775A2D90A";
   constant CPIX_NORMAL_INIT_1C_BIT_13_C : bit_vector(255 downto 0) := x"875F5BE6CC7221DF3078795AD62661B388B665CFB07BDBC416660BCFAA1D63D4";
   constant CPIX_NORMAL_INIT_1C_BIT_14_C : bit_vector(255 downto 0) := x"BB647FE4F05AC85A20FB05135F26D084578AB031FB65DEA45DA9C8B9760DFDDD";
   constant CPIX_NORMAL_INIT_1D_BIT_00_C : bit_vector(255 downto 0) := x"E5511D84245C8EC052ECFB24F8F28D31A058F0704A33D84D5F9772ACC75C6CE2";
   constant CPIX_NORMAL_INIT_1D_BIT_01_C : bit_vector(255 downto 0) := x"40ADB75E64028511C1E314CB1C087C5C29E872BE516AF39975B6D5613BDC200F";
   constant CPIX_NORMAL_INIT_1D_BIT_02_C : bit_vector(255 downto 0) := x"79833D3080F7A439AED43E3F7FD53C16669F9F0E2FCB433DF69C52C998D76CEC";
   constant CPIX_NORMAL_INIT_1D_BIT_03_C : bit_vector(255 downto 0) := x"BB7FA4921BB6AC4514D158272B952AE2CF2D70F914D05571F4D888B9E4FA1A65";
   constant CPIX_NORMAL_INIT_1D_BIT_04_C : bit_vector(255 downto 0) := x"3161AC94050E0E6ADC060BCED9800F1BD2FA6E8C48614CE42F97EB46132CEC68";
   constant CPIX_NORMAL_INIT_1D_BIT_05_C : bit_vector(255 downto 0) := x"10CD24A7C50D75515DC108C8D58072E87AC1BF621C30F6A95C92DF5D16053BBA";
   constant CPIX_NORMAL_INIT_1D_BIT_06_C : bit_vector(255 downto 0) := x"0725EEC23C56AEF4DD8256B5120232A75031A79956C80D5536F2714B7A286CFD";
   constant CPIX_NORMAL_INIT_1D_BIT_07_C : bit_vector(255 downto 0) := x"30330670E151ABB77EE9C68C82464D83F945FBA03CDD31466C3A91A712878569";
   constant CPIX_NORMAL_INIT_1D_BIT_08_C : bit_vector(255 downto 0) := x"E1A4D63FB74CD6BB733E63423DA56E9D23D1D5E1D79AFD9A48CF079C3CA48AF9";
   constant CPIX_NORMAL_INIT_1D_BIT_09_C : bit_vector(255 downto 0) := x"B4306A4FF2A61EE295BC2D79241EAC65A1B8BF9D1079776572E90C31486171B2";
   constant CPIX_NORMAL_INIT_1D_BIT_10_C : bit_vector(255 downto 0) := x"D081C14087D8A67D02B837349B64D971313A48BE8BAC2565ED4239A28E1B786D";
   constant CPIX_NORMAL_INIT_1D_BIT_11_C : bit_vector(255 downto 0) := x"85F50E57222FCF07883994D00525948460A0BD523063347480FADCC655AA175B";
   constant CPIX_NORMAL_INIT_1D_BIT_12_C : bit_vector(255 downto 0) := x"30CAFA7F3535601BC0F78B87EC993AECB7EAECDB8217CF5E0A21CA4DB40FC033";
   constant CPIX_NORMAL_INIT_1D_BIT_13_C : bit_vector(255 downto 0) := x"2BB8EDAFB0FD9B691BA5CE4769F9CA5E417DFBB0880730E95044364BCED6901D";
   constant CPIX_NORMAL_INIT_1D_BIT_14_C : bit_vector(255 downto 0) := x"3905A60F1E674DBDDFC69D6C2CDB035FBC78DF464D698549F5D7D98AF5D008A4";
   constant CPIX_NORMAL_INIT_1E_BIT_00_C : bit_vector(255 downto 0) := x"C4DDAA3AE1ADF6B1EA0EA5288F7FCDB5D377EE3B782A06C384A0D329CCDCC6FC";
   constant CPIX_NORMAL_INIT_1E_BIT_01_C : bit_vector(255 downto 0) := x"45E20E96E27DEED9EC60AC91A389E5D94DCAE927A764B519034484D14462A7D2";
   constant CPIX_NORMAL_INIT_1E_BIT_02_C : bit_vector(255 downto 0) := x"7FEB894281CC11BE006D1BAD8A96BC8FB0236F22F126D86EAC9796DDB6ECCC17";
   constant CPIX_NORMAL_INIT_1E_BIT_03_C : bit_vector(255 downto 0) := x"C88697713886A7CAAC2CF4C7F36F6205188F2217740CDB455F39E1DD2B9F5578";
   constant CPIX_NORMAL_INIT_1E_BIT_04_C : bit_vector(255 downto 0) := x"0BFA54E4062F1F3334CF3385F2DA31AD32BC40F353DA98720DB7AD6D1FE9B678";
   constant CPIX_NORMAL_INIT_1E_BIT_05_C : bit_vector(255 downto 0) := x"834144FB53E309A6DB9DE4238C45936F4C9F1FD011570D7A4C1FA6487C0FCA34";
   constant CPIX_NORMAL_INIT_1E_BIT_06_C : bit_vector(255 downto 0) := x"EE65FC2A99D33DCD82623E362E5A14F61950A5E173414377159C6AD9A5C501C3";
   constant CPIX_NORMAL_INIT_1E_BIT_07_C : bit_vector(255 downto 0) := x"D1B417085DEF695DC5582C5955FEA6BB11690A963EAC3AD15BC768CDBAA7BB1E";
   constant CPIX_NORMAL_INIT_1E_BIT_08_C : bit_vector(255 downto 0) := x"628ED2F46443A8B792314E5A308B882D1DEF2E207C73E9F9395CF083912F618F";
   constant CPIX_NORMAL_INIT_1E_BIT_09_C : bit_vector(255 downto 0) := x"3843FEF349A1308C39B326AFF641A0586B8056DE11835EE10AD1538CD49CCC9E";
   constant CPIX_NORMAL_INIT_1E_BIT_10_C : bit_vector(255 downto 0) := x"A315860E578200751F996B55531FFBF225AE3C820451DC8A41A84D0855E1188B";
   constant CPIX_NORMAL_INIT_1E_BIT_11_C : bit_vector(255 downto 0) := x"E45E2016122B1B198F4AEB2ED4753225A715E00B7EBF0D7C1F60683C73A6FE56";
   constant CPIX_NORMAL_INIT_1E_BIT_12_C : bit_vector(255 downto 0) := x"CA2813091CB71D050EB5B8ED9E8BDF8032B7D35FBAF999E55A8D1EE144F95034";
   constant CPIX_NORMAL_INIT_1E_BIT_13_C : bit_vector(255 downto 0) := x"C1B37503966AC24F123693A1AA4213130AEEC0BBFDE95639D9C792D722ED080F";
   constant CPIX_NORMAL_INIT_1E_BIT_14_C : bit_vector(255 downto 0) := x"588A95F6B3DA20B920DBB836A42BBB0E2139A7F99B5C7D402308E4FA2418B996";
   constant CPIX_NORMAL_INIT_1F_BIT_00_C : bit_vector(255 downto 0) := x"CFA1FCE35944F24ADDDE7E3FED02115A25188A8A2C8E653C4B27ED9D5185CB9A";
   constant CPIX_NORMAL_INIT_1F_BIT_01_C : bit_vector(255 downto 0) := x"5390EE0C558AFBA531A88626636BD2F9BE1876B061B417195935CF9DD2143429";
   constant CPIX_NORMAL_INIT_1F_BIT_02_C : bit_vector(255 downto 0) := x"B66E2DD7AC132C31CD4A22B79298F817FD3D0583A168929BB51F99AA36C895DC";
   constant CPIX_NORMAL_INIT_1F_BIT_03_C : bit_vector(255 downto 0) := x"FFBFF963B2F10FE74CEC7D95757BCD1CC360E4F960F63A40AE971442BC2D8449";
   constant CPIX_NORMAL_INIT_1F_BIT_04_C : bit_vector(255 downto 0) := x"11CE216A096855E510EE8170450F708DB80ED2CE07AC34FCB8FE9D4AE26A08C7";
   constant CPIX_NORMAL_INIT_1F_BIT_05_C : bit_vector(255 downto 0) := x"56F91E720C055B93126449F122BE8D43325A1F876D133339C088741EA3585230";
   constant CPIX_NORMAL_INIT_1F_BIT_06_C : bit_vector(255 downto 0) := x"1C892FC75E29562309B8961720DB3FC19CA08E461807230F16787B77AD3EB36C";
   constant CPIX_NORMAL_INIT_1F_BIT_07_C : bit_vector(255 downto 0) := x"162938CB10E7C860AAC505DF74276453D5EB1FCAA722F75C2B487DAF0DDD44C3";
   constant CPIX_NORMAL_INIT_1F_BIT_08_C : bit_vector(255 downto 0) := x"3674299F56BC24F52868A01032E7EF5F3F7724DF0F0AC893B4E8D65BAB06AC99";
   constant CPIX_NORMAL_INIT_1F_BIT_09_C : bit_vector(255 downto 0) := x"10A5BB1E50F32EC17BB1F2768C9CC6B63EEB6722992B48CEA8400D7EDD958054";
   constant CPIX_NORMAL_INIT_1F_BIT_10_C : bit_vector(255 downto 0) := x"018F3B724DC435B7627716968242DE2F215B58E22F20E534A1A0BED598E2377B";
   constant CPIX_NORMAL_INIT_1F_BIT_11_C : bit_vector(255 downto 0) := x"10C743D6414E61F055A93C609CB96F4B8CA9D5F41E880BA090293BF90236BF14";
   constant CPIX_NORMAL_INIT_1F_BIT_12_C : bit_vector(255 downto 0) := x"128209D908721D726776052CA17443FD1E1AC30922E94E1C0322FB3C8F6E800B";
   constant CPIX_NORMAL_INIT_1F_BIT_13_C : bit_vector(255 downto 0) := x"106328DC34087728379297D002ACAF4CA505106C275FF39E125F95B193E33DBA";
   constant CPIX_NORMAL_INIT_1F_BIT_14_C : bit_vector(255 downto 0) := x"02411A89C188BC4A354B30472455C4D36CC2DE075B293AEEC77F283BD4C2F4BB";
   constant CPIX_NORMAL_INIT_20_BIT_00_C : bit_vector(255 downto 0) := x"74AA3C8EC1969FEAFE8874662B5329189DEA15E756EA049B4081D9F647682A93";
   constant CPIX_NORMAL_INIT_20_BIT_01_C : bit_vector(255 downto 0) := x"2E5910845FD033DC29DEEC51BC972A7F305BC858236F4006DE33A5FD1DF00D6A";
   constant CPIX_NORMAL_INIT_20_BIT_02_C : bit_vector(255 downto 0) := x"7485ECE03F1279F15F9E9D57ACFB20E3B82C25D1C98B8E5B9528DC17F66FAFDB";
   constant CPIX_NORMAL_INIT_20_BIT_03_C : bit_vector(255 downto 0) := x"1CEF6613EC0DCD59B290A0BC88A79A32E2F952C058A9350DB96EB8FA43ECA47B";
   constant CPIX_NORMAL_INIT_20_BIT_04_C : bit_vector(255 downto 0) := x"4935C88338AD9645C027BF01183C3CA9A368B4A33B4FCB0CF23E34C7CF15CB69";
   constant CPIX_NORMAL_INIT_20_BIT_05_C : bit_vector(255 downto 0) := x"68CDF565207A52725E9B273B36E40B91E546D68B5909051DFADE0093D7339D97";
   constant CPIX_NORMAL_INIT_20_BIT_06_C : bit_vector(255 downto 0) := x"905EB9A276C24C856BB600A8F0C06903B0CDF8A167DEFFD2C1317133577FF43B";
   constant CPIX_NORMAL_INIT_20_BIT_07_C : bit_vector(255 downto 0) := x"AB1A7AFA8F7D5299FDB27E6749A617F305DE7ACC3AA0FC9499A8C6694AD0D57F";
   constant CPIX_NORMAL_INIT_20_BIT_08_C : bit_vector(255 downto 0) := x"CDC75FA8457196673A21ED73D6F150FB7EF8879C7C3986DBD001FEE7C9F8FFCF";
   constant CPIX_NORMAL_INIT_20_BIT_09_C : bit_vector(255 downto 0) := x"54EF4960C0914D6213169F1B25EE8F05550C9DF3BB813E8173C78F18C7BCFE63";
   constant CPIX_NORMAL_INIT_20_BIT_10_C : bit_vector(255 downto 0) := x"6A1D0A0EAEC7FA3EA11815EA021B555966C2EACC15FE5B41CE0E9C85F97AF631";
   constant CPIX_NORMAL_INIT_20_BIT_11_C : bit_vector(255 downto 0) := x"CE0032768A66FC9D3050DE46DFD8C42C11CB319E0E0F7373A1CAF47BECD02FA3";
   constant CPIX_NORMAL_INIT_20_BIT_12_C : bit_vector(255 downto 0) := x"9036386A150F596C99EE8AF853E3AE6616359A743C31FA44EE58ABC156DA3307";
   constant CPIX_NORMAL_INIT_20_BIT_13_C : bit_vector(255 downto 0) := x"A72A8CDF54262146BDA71CF4F17E87D468D2EFBC255A23B6678F7854004E5BE3";
   constant CPIX_NORMAL_INIT_20_BIT_14_C : bit_vector(255 downto 0) := x"95CB439744175EB060D97F183A8A6370D52F5D76857B56FD64A287A8A19B11A5";
   constant CPIX_NORMAL_INIT_21_BIT_00_C : bit_vector(255 downto 0) := x"1DF5EE672896072940A92A62694C3D6E65B9FBECA8A5632FB4E274A4AFF4F530";
   constant CPIX_NORMAL_INIT_21_BIT_01_C : bit_vector(255 downto 0) := x"6B953390C7F3FD3750BD990B32840D412C49C0073CC469BF052BAFDD5DB572F2";
   constant CPIX_NORMAL_INIT_21_BIT_02_C : bit_vector(255 downto 0) := x"754042E9EB025E4D64F49D37F147FEAC522EF0ED0D98F14D94F8AD8837651516";
   constant CPIX_NORMAL_INIT_21_BIT_03_C : bit_vector(255 downto 0) := x"FE0358466BCC9C2A4873585907DAC36D93341D49CDF21B0B554BF77F3B04751C";
   constant CPIX_NORMAL_INIT_21_BIT_04_C : bit_vector(255 downto 0) := x"9FFEEBE75EC3C274037A2F296F172638CE0EC3B5FFFC44092A2D972C07ABFC8E";
   constant CPIX_NORMAL_INIT_21_BIT_05_C : bit_vector(255 downto 0) := x"969E09DEEF15D3DE97C558077D68528EF71E5ACE1A32A0321FCE2DDB0F52AE1F";
   constant CPIX_NORMAL_INIT_21_BIT_06_C : bit_vector(255 downto 0) := x"BE1B524C4A67495F47F2D357ECA8616AE535400273EB5FF30DABD140A82D21E8";
   constant CPIX_NORMAL_INIT_21_BIT_07_C : bit_vector(255 downto 0) := x"D0DE7FE54629C9AAD62320273782F1ABEC64C4D953C4A31CB620FE8ADBEBFBDC";
   constant CPIX_NORMAL_INIT_21_BIT_08_C : bit_vector(255 downto 0) := x"796D87DB3B3DA4569D1C134B831BA1AC2077D2220480D806BFD92AAE108FB39F";
   constant CPIX_NORMAL_INIT_21_BIT_09_C : bit_vector(255 downto 0) := x"52B415074CE8725BC168E7E102EE7B59DD9E8A8BDB3C305472A1F27772D1080C";
   constant CPIX_NORMAL_INIT_21_BIT_10_C : bit_vector(255 downto 0) := x"91814A9D38E36A54F442D83C39E89F5A06D2670AD1A661697B2566F70E08822A";
   constant CPIX_NORMAL_INIT_21_BIT_11_C : bit_vector(255 downto 0) := x"3BACBC74280B0371078B265A44CA7648B417D5773553F5A2B766379A4D4D0649";
   constant CPIX_NORMAL_INIT_21_BIT_12_C : bit_vector(255 downto 0) := x"55F7C66AD3D63DE110B5863B0E9DD7D705B73079E513CF47279932C7F5185222";
   constant CPIX_NORMAL_INIT_21_BIT_13_C : bit_vector(255 downto 0) := x"637930F3F3959C6688BE0A8D1CF2F3F01FB8B9F35A843DCE4292E74F96B0BDBD";
   constant CPIX_NORMAL_INIT_21_BIT_14_C : bit_vector(255 downto 0) := x"783DBBEE57B4388FEF13198BB0B9BCDBA56399E7C8BB937A4728894EC691F9C7";
   constant CPIX_NORMAL_INIT_22_BIT_00_C : bit_vector(255 downto 0) := x"0EFA510DA504CF21E6E74E21AF3C4358C829A7FFBB3D3148DBD4C3F01BD0D9B2";
   constant CPIX_NORMAL_INIT_22_BIT_01_C : bit_vector(255 downto 0) := x"49CD707723821FCC7638155F932AB2670D905B075A244E1FC28D9E1E0C9C99E5";
   constant CPIX_NORMAL_INIT_22_BIT_02_C : bit_vector(255 downto 0) := x"E68FA36B86402415DB656AD8C2FA9A608C26D9DBCDCB7895DD92399BAE03F544";
   constant CPIX_NORMAL_INIT_22_BIT_03_C : bit_vector(255 downto 0) := x"10AE609D6AAB29FF244AEA853E8308D1AE8EF121E4F33772E41AC110995E41FB";
   constant CPIX_NORMAL_INIT_22_BIT_04_C : bit_vector(255 downto 0) := x"1A488FC96A654D1B524A1B9B4E60EA5D638BB6DEE1E1F4BFB1CFDCCF05BD62F9";
   constant CPIX_NORMAL_INIT_22_BIT_05_C : bit_vector(255 downto 0) := x"5A363F0E64A120943996B6455C2F3E88B479EA23E249FF0547B343A3D3CDEC38";
   constant CPIX_NORMAL_INIT_22_BIT_06_C : bit_vector(255 downto 0) := x"EBB3AE12B939063777CDEFDE1B020A23DC43839B392F58B12D192C6ED32BC4A3";
   constant CPIX_NORMAL_INIT_22_BIT_07_C : bit_vector(255 downto 0) := x"9157A0D41038A8D7780FF9D845208B5F232E56C876C5F14D1CFC2DDDB157B0CD";
   constant CPIX_NORMAL_INIT_22_BIT_08_C : bit_vector(255 downto 0) := x"D861CBB4281B171F16F22D0F258A203D00AC25CFFDF007DAC2AD37DEEF0F41F3";
   constant CPIX_NORMAL_INIT_22_BIT_09_C : bit_vector(255 downto 0) := x"D01D3996397E83C669682C2F6BBBD6E30AB2AD1E8E2F963D22ADAE7C3BE18686";
   constant CPIX_NORMAL_INIT_22_BIT_10_C : bit_vector(255 downto 0) := x"648A580B53BB5D33770CBA3E167EFF4FD755609EDE2E7B36AEEBEF6D4753DF6A";
   constant CPIX_NORMAL_INIT_22_BIT_11_C : bit_vector(255 downto 0) := x"7EFF2237750D308C896B09489E0DDD6A1D77D9E0A58546B25078BF0DAF0713EC";
   constant CPIX_NORMAL_INIT_22_BIT_12_C : bit_vector(255 downto 0) := x"E934676AAE3D8103E3B6EC7A611ED5DB8F47FAE24151E61B62DA671F464A7C0A";
   constant CPIX_NORMAL_INIT_22_BIT_13_C : bit_vector(255 downto 0) := x"29D309DBB7F970441E858E85C8D0FEF1B6B2C051F4C39E44F7F9600D8C95C26A";
   constant CPIX_NORMAL_INIT_22_BIT_14_C : bit_vector(255 downto 0) := x"0248CEDCC8C73D7E45051470BDD33CFBB707CF77041FE31603A8D12ED73C8EB6";
   constant CPIX_NORMAL_INIT_23_BIT_00_C : bit_vector(255 downto 0) := x"6C8ACB3CCD3308DDFD5BF31617D958CADAED054C5234AF5A49360B6AD8370771";
   constant CPIX_NORMAL_INIT_23_BIT_01_C : bit_vector(255 downto 0) := x"354B96EB48C4AFA536F43AA0465DDE86D5FABF76C0F64F32AF2F48FBB890A05D";
   constant CPIX_NORMAL_INIT_23_BIT_02_C : bit_vector(255 downto 0) := x"A9B2CCA71CDADA94BB46051208A8D7127633E74AEE4BAA924AAD091B0922BECB";
   constant CPIX_NORMAL_INIT_23_BIT_03_C : bit_vector(255 downto 0) := x"F2864A776BCCF818675D8114DAE5663E4A583532CA61B992287DEB06B5E3DB11";
   constant CPIX_NORMAL_INIT_23_BIT_04_C : bit_vector(255 downto 0) := x"70C6307AC7AC155A2437E1E842F257DA1BB9AA8D5235D9EFB96B6D2D6FC7C07A";
   constant CPIX_NORMAL_INIT_23_BIT_05_C : bit_vector(255 downto 0) := x"930FF6389D1365763006B36B48EE426C919AD2C48FD91AAD15C0D6402995523D";
   constant CPIX_NORMAL_INIT_23_BIT_06_C : bit_vector(255 downto 0) := x"3B34379694FD0B31966B29D8F6D1CE781B623CE291338109724FC6F3919845EF";
   constant CPIX_NORMAL_INIT_23_BIT_07_C : bit_vector(255 downto 0) := x"94957E9124073ADF63AD205C89C14182C3AB61BE59390828E36F25CF2A81ECA2";
   constant CPIX_NORMAL_INIT_23_BIT_08_C : bit_vector(255 downto 0) := x"980FDD3CE5B464053BF28D62EA5A86C50BFA900590FE1E320E2FB97C8A90C44D";
   constant CPIX_NORMAL_INIT_23_BIT_09_C : bit_vector(255 downto 0) := x"36B3F5107078B6A13F042281E08E52A2615D6274C1BF2A03F8BF1D9E38A3311F";
   constant CPIX_NORMAL_INIT_23_BIT_10_C : bit_vector(255 downto 0) := x"71FF5827BCAF51010AA8585C252FF3232A6E6F9C3D683DF4154F6886D419B778";
   constant CPIX_NORMAL_INIT_23_BIT_11_C : bit_vector(255 downto 0) := x"74030A2E5EF29C8F3F00145777E1FB754C94CDCFBF6F6FFFAF1F6676ECE63E84";
   constant CPIX_NORMAL_INIT_23_BIT_12_C : bit_vector(255 downto 0) := x"C5C2EAEDA48EF8A07172DFA50C5A7295DC0F8D1FA750EFDD7D9BF070B50F7AB7";
   constant CPIX_NORMAL_INIT_23_BIT_13_C : bit_vector(255 downto 0) := x"42EA0FCD5FEFD27992B3243CF51D56FA9D6F370B0FD977DC064856F416A5306B";
   constant CPIX_NORMAL_INIT_23_BIT_14_C : bit_vector(255 downto 0) := x"A1517BD55C5728913CC73050A55CCA081A0E4F6075DBB5F4FF8A6FA79DD33C63";
   constant CPIX_NORMAL_INIT_24_BIT_00_C : bit_vector(255 downto 0) := x"C826E76655DA7CB97420EB758BD33CA99B8674893D15C756C9CEDCB7A863A2E4";
   constant CPIX_NORMAL_INIT_24_BIT_01_C : bit_vector(255 downto 0) := x"D6D13B6E16F0C1D1390974AFCC3D11E316D2FCA6DC7503199B29322BDDDB10DA";
   constant CPIX_NORMAL_INIT_24_BIT_02_C : bit_vector(255 downto 0) := x"CABC2890D58136E14E24A9FD4D7C1ADFC905033805DB9303F5F93EB6F12EB5E1";
   constant CPIX_NORMAL_INIT_24_BIT_03_C : bit_vector(255 downto 0) := x"F237A5CD0960F4F2B52C1CF88C7D499B718F991E483D444608A7B9CE81AD10B9";
   constant CPIX_NORMAL_INIT_24_BIT_04_C : bit_vector(255 downto 0) := x"E679B14FE4F2AF549E72F0D89AB44C50584BA945A9EBF150FE4FD02B93488E7A";
   constant CPIX_NORMAL_INIT_24_BIT_05_C : bit_vector(255 downto 0) := x"25BD629C45D357C234ABCC0B2F6A7ECCE5766A22F0673AF8DB92EDDD86F270FD";
   constant CPIX_NORMAL_INIT_24_BIT_06_C : bit_vector(255 downto 0) := x"22064D4A607D24E2ADAD9E41D901C422B2CAD4F1F3BE741DEDF11F40DCC10F3D";
   constant CPIX_NORMAL_INIT_24_BIT_07_C : bit_vector(255 downto 0) := x"347DC09B7E09651591E064741000843C2781D0D94143E80469DD0ABE7A776809";
   constant CPIX_NORMAL_INIT_24_BIT_08_C : bit_vector(255 downto 0) := x"FFE4D7F48A03537E37329BBCAFEF6A1B40DEC7C827D413BD393C71B76399A333";
   constant CPIX_NORMAL_INIT_24_BIT_09_C : bit_vector(255 downto 0) := x"B3992B34BD27BBA832563EDFA6FFEFC7C2A72755171FDEAB932E78B841F61AEB";
   constant CPIX_NORMAL_INIT_24_BIT_10_C : bit_vector(255 downto 0) := x"E77078FC9E8C928B317CC3B28B3F57DB5487E0525DBF9FEF2643F4BBBF1CE6C6";
   constant CPIX_NORMAL_INIT_24_BIT_11_C : bit_vector(255 downto 0) := x"CBC7ADD8DEF2DA46FA25C23BCFBF73D37D9A1FF6F049432E86F655F2BC385F53";
   constant CPIX_NORMAL_INIT_24_BIT_12_C : bit_vector(255 downto 0) := x"D609CDBACBCA37C0A2902F3C9EAF727764665A4739D5F3FD7C3B47B3546FA2AF";
   constant CPIX_NORMAL_INIT_24_BIT_13_C : bit_vector(255 downto 0) := x"A71E19717876838DFE382259C6AFE747EEC37AA958A2C683996699F8D54667C7";
   constant CPIX_NORMAL_INIT_24_BIT_14_C : bit_vector(255 downto 0) := x"13EB506BCC1DCED2A9B1AA10D32F432E2442E4F5A505F79B39D15799762E5664";
   constant CPIX_NORMAL_INIT_25_BIT_00_C : bit_vector(255 downto 0) := x"FF5914A56E09070F4F8F5913BA0F8B0EB471E4A719FE343D9FA9D9991AE4FEE8";
   constant CPIX_NORMAL_INIT_25_BIT_01_C : bit_vector(255 downto 0) := x"AFD003DAEC813AED526A596784AFB6A4C092FEC46D68A044C1F05ADC15423992";
   constant CPIX_NORMAL_INIT_25_BIT_02_C : bit_vector(255 downto 0) := x"F954532354F8E3AA65D5E1F1464F00A799D2F86601FF779D2D8480DD99D1E610";
   constant CPIX_NORMAL_INIT_25_BIT_03_C : bit_vector(255 downto 0) := x"BAC65E06C34941A6F9A96C05A352FC9C72457B93EDAE541F0469C4A46406DD63";
   constant CPIX_NORMAL_INIT_25_BIT_04_C : bit_vector(255 downto 0) := x"43D0C96713DDF2214846E18AD9353BA9BEF3B3365FBC184094F0CAF1D17D8400";
   constant CPIX_NORMAL_INIT_25_BIT_05_C : bit_vector(255 downto 0) := x"6C71B7C700DDAC34C381FCB02AE9AB4367DF2190AFC75C71325AAD07C1414377";
   constant CPIX_NORMAL_INIT_25_BIT_06_C : bit_vector(255 downto 0) := x"821D1E98ABE885DA275CC9649F43E1EA0F81B10A072AAB95902E440DF2EC6407";
   constant CPIX_NORMAL_INIT_25_BIT_07_C : bit_vector(255 downto 0) := x"12E0508EA43ACCBFA68265DCED692091E89E5BE95822D9D4D58277FAE8F20DD5";
   constant CPIX_NORMAL_INIT_25_BIT_08_C : bit_vector(255 downto 0) := x"6D89E36A6D0BBA0E1439A8BF3C85C6597EA81DEA0BFDCF1EBB6037F786D7C13C";
   constant CPIX_NORMAL_INIT_25_BIT_09_C : bit_vector(255 downto 0) := x"B19CBA92F4A0B284750FD3CEC43FE3F538E1B262B7EFDA74678F94AA8B8E562A";
   constant CPIX_NORMAL_INIT_25_BIT_10_C : bit_vector(255 downto 0) := x"B80DAB4E208548DE04EF2FCF8FEF3864C6632435618D3AD236894FBA2D6CF251";
   constant CPIX_NORMAL_INIT_25_BIT_11_C : bit_vector(255 downto 0) := x"AE7A9B22EAD9EE706931EECC646684AE4ADB5D60BDF162B4A9B046BB3684EACE";
   constant CPIX_NORMAL_INIT_25_BIT_12_C : bit_vector(255 downto 0) := x"3FD56258F9F587656BA024A6BD34C1A92C443B5DC3A6C34A3C618AB61F363828";
   constant CPIX_NORMAL_INIT_25_BIT_13_C : bit_vector(255 downto 0) := x"360E8E8B0AAA56ADB1415F8F53D19070A5A8A359B074AAD059F21DA2769899BE";
   constant CPIX_NORMAL_INIT_25_BIT_14_C : bit_vector(255 downto 0) := x"82D08780FAE1B946ABA40B2E08F17C563250FAC4BF152E6DA92D116EE4FD14FC";
   constant CPIX_NORMAL_INIT_26_BIT_00_C : bit_vector(255 downto 0) := x"238DFF643F49B7518460726DC8BE38DA2FD959CCF809DA9AD4BEC5399D9E92CD";
   constant CPIX_NORMAL_INIT_26_BIT_01_C : bit_vector(255 downto 0) := x"02A1768B028639B91ECF7443B8BF153EC032849005158F40BBB5312E945E8EDA";
   constant CPIX_NORMAL_INIT_26_BIT_02_C : bit_vector(255 downto 0) := x"6A54BD759C58D3301872578E9779B312AA135510E6DD93C21101901F8771A990";
   constant CPIX_NORMAL_INIT_26_BIT_03_C : bit_vector(255 downto 0) := x"CCB7D197AB6B7511523F87A1B085F5A5339B19398C484C19186D2566C52C56D7";
   constant CPIX_NORMAL_INIT_26_BIT_04_C : bit_vector(255 downto 0) := x"B326AF59148A35F357B7A2AB4C987F588BE9B04F075142AE4FDC5E8A3CCA41ED";
   constant CPIX_NORMAL_INIT_26_BIT_05_C : bit_vector(255 downto 0) := x"74A7F5AC912E94BBF29ED917392CB21340A6F3132939BBA38BE584B025B8664C";
   constant CPIX_NORMAL_INIT_26_BIT_06_C : bit_vector(255 downto 0) := x"F9B75B8510F57521B0D2EE92AB9F692BCCBD5E54CC24141D4FED9294D03D7E8D";
   constant CPIX_NORMAL_INIT_26_BIT_07_C : bit_vector(255 downto 0) := x"844F8E5AA392EF08D5E07DECBB9C3007745E87CDF9800D26B86FCD56C893DC46";
   constant CPIX_NORMAL_INIT_26_BIT_08_C : bit_vector(255 downto 0) := x"1A7005C163EC6FB42934BD3C2960DA8BD0EEA5AE05C7E203957A8A4B16CE3FAC";
   constant CPIX_NORMAL_INIT_26_BIT_09_C : bit_vector(255 downto 0) := x"FF6C3ED79B4E7067E45D5FC9D416870FC3E563163F845B7B068C8B5DB379D1F5";
   constant CPIX_NORMAL_INIT_26_BIT_10_C : bit_vector(255 downto 0) := x"5B91095BDF5F270137001CE47F073D45F2ACE916A485DEA95AC8F12DEEBD66D7";
   constant CPIX_NORMAL_INIT_26_BIT_11_C : bit_vector(255 downto 0) := x"5AFB893F1FF3F288664F6AD694C1B67D53FA852F0B18DBC0FDF70DC4F9328B41";
   constant CPIX_NORMAL_INIT_26_BIT_12_C : bit_vector(255 downto 0) := x"0E1E55C8069C4F1B9FDADC158E8827E4AC2CFA8E389F8F02D3B7A861E1CCF9D5";
   constant CPIX_NORMAL_INIT_26_BIT_13_C : bit_vector(255 downto 0) := x"3D2A5BBFD3503D75DCB7A6729D8766B4D200F12DFD41424EDAA00DF11796A44A";
   constant CPIX_NORMAL_INIT_26_BIT_14_C : bit_vector(255 downto 0) := x"426F240C62D6DC24DC0C6CFF2E7B3D4AD2A321B8EAFBAF182243B50ABCC81238";
   constant CPIX_NORMAL_INIT_27_BIT_00_C : bit_vector(255 downto 0) := x"59C8EB4E600657D6325B0477F3810D227C208CA72A39F860C3982082AE8109AE";
   constant CPIX_NORMAL_INIT_27_BIT_01_C : bit_vector(255 downto 0) := x"1F323FA455900856BDCCFCA8BAB0BCF9E1F8A675B530121EABE2525311974283";
   constant CPIX_NORMAL_INIT_27_BIT_02_C : bit_vector(255 downto 0) := x"98017C0FA0DBF4D86982E1812E78877A3FCB8D8F8967BBAE4B9FF796128207B9";
   constant CPIX_NORMAL_INIT_27_BIT_03_C : bit_vector(255 downto 0) := x"E5B533F243B838C12604E951B9BD7306D3293D75DA8FB1274F7E6C24B7C2E0B6";
   constant CPIX_NORMAL_INIT_27_BIT_04_C : bit_vector(255 downto 0) := x"C44DB65988DAAC41481F7DAD8BDA75DAD34880C2201064C6385AF8ADD747B62E";
   constant CPIX_NORMAL_INIT_27_BIT_05_C : bit_vector(255 downto 0) := x"BA1FB725ADEF0A2A53D4911D36E630929057D0C89CA9AF986A1DAD9642BBB5EC";
   constant CPIX_NORMAL_INIT_27_BIT_06_C : bit_vector(255 downto 0) := x"95995B3D8015AF6C18FD0A2AE5D7E35550A2CB89B787AD83B9F78D01FB8893E8";
   constant CPIX_NORMAL_INIT_27_BIT_07_C : bit_vector(255 downto 0) := x"99900793DC4E4D71ECD763E3D28BD19EB2779005DCBC2D95622D71AEC3096F33";
   constant CPIX_NORMAL_INIT_27_BIT_08_C : bit_vector(255 downto 0) := x"A7A30297F3438B430A13B291D0B7E9D54BCBE4D37DEE1683830A76BF59B3A090";
   constant CPIX_NORMAL_INIT_27_BIT_09_C : bit_vector(255 downto 0) := x"9EB1FA2294D006F29B58F1924AD93CA2A188E7216FBD931E24E4739608AB6431";
   constant CPIX_NORMAL_INIT_27_BIT_10_C : bit_vector(255 downto 0) := x"5E4F3A0978464B8F70C3F7FE483844D994632ECFE2454C39DBB6E7DEBAE67489";
   constant CPIX_NORMAL_INIT_27_BIT_11_C : bit_vector(255 downto 0) := x"9646D8B51E849F2E229F44B971B6C2CA73153A580E9A28CF2212FD8FDEB9DCD8";
   constant CPIX_NORMAL_INIT_27_BIT_12_C : bit_vector(255 downto 0) := x"872E6467A5124E410DBD399CBFBD993A8BF33538C3361193D2C4E6CF9F1DCBCC";
   constant CPIX_NORMAL_INIT_27_BIT_13_C : bit_vector(255 downto 0) := x"928CEE04587EBFDE7D81AD0F03DBDB1165BDD1727E19892B7C27AE8725BC8536";
   constant CPIX_NORMAL_INIT_27_BIT_14_C : bit_vector(255 downto 0) := x"1948D93309D8738B8EE33A1C77EC422ED197CC37AC55FCE0CCA237C8CBD8D39F";
   constant CPIX_NORMAL_INIT_28_BIT_00_C : bit_vector(255 downto 0) := x"0673FEF894A664B72D45116617FCE6EEF125104C7C15886E886C8876CD831E43";
   constant CPIX_NORMAL_INIT_28_BIT_01_C : bit_vector(255 downto 0) := x"26FA57C711D9AC5CA4B35036927CE5D28180427AEE78A805C7119C4C4DAF481B";
   constant CPIX_NORMAL_INIT_28_BIT_02_C : bit_vector(255 downto 0) := x"475091C9A5CBBB15B1B0821E9D270ACE40C96DA267150CDB57FE737DCAFC838C";
   constant CPIX_NORMAL_INIT_28_BIT_03_C : bit_vector(255 downto 0) := x"851A67532FD79CCB23A701859D1A262598C87B478B7DD7CFD407B2567031CA4B";
   constant CPIX_NORMAL_INIT_28_BIT_04_C : bit_vector(255 downto 0) := x"8E5E356FF07C5D52A5B78F07CA5BD973E512257005F11C5935990DED09F4A97D";
   constant CPIX_NORMAL_INIT_28_BIT_05_C : bit_vector(255 downto 0) := x"DEE68C41E839C07B8CB2E99C311D75D2A67ED9C8E8B2C762192AB7C349F7A3F7";
   constant CPIX_NORMAL_INIT_28_BIT_06_C : bit_vector(255 downto 0) := x"EAB796F3C8F593E57253D6C597DB70D1B8176F0470CF5C14AC8160C5994E7FFB";
   constant CPIX_NORMAL_INIT_28_BIT_07_C : bit_vector(255 downto 0) := x"BB1B521556F05510F2A39E43489DA7F9AD1491CD03C688DE6A7BE90F688AC12F";
   constant CPIX_NORMAL_INIT_28_BIT_08_C : bit_vector(255 downto 0) := x"9E61E42069AA1E21963FA54305E61E57D7F2ED743808F09F5C7997BBA6B3996D";
   constant CPIX_NORMAL_INIT_28_BIT_09_C : bit_vector(255 downto 0) := x"BEA9C1087271BE9FBEE44179261B12D0AD0B450FE1EA9BB09434EF45CFD9D669";
   constant CPIX_NORMAL_INIT_28_BIT_10_C : bit_vector(255 downto 0) := x"F99D0A5D06CED0BE09FFCAADF28E157CD3928ACE24C5D300301A6C3F00ED09EB";
   constant CPIX_NORMAL_INIT_28_BIT_11_C : bit_vector(255 downto 0) := x"90A9CBDF25D77208B3D8549CFC52AD5CCA175208BFFCCE510A0BA8E0DE1F4B25";
   constant CPIX_NORMAL_INIT_28_BIT_12_C : bit_vector(255 downto 0) := x"4108ED2B9767FADB6435626F58732708F0EDB33F7B7579E8A8DCC2D0BAB825AD";
   constant CPIX_NORMAL_INIT_28_BIT_13_C : bit_vector(255 downto 0) := x"05DBB2FADD7E0A9977F8912BA398F1307BF821AEEF8C25AF4384DAE626665A0D";
   constant CPIX_NORMAL_INIT_28_BIT_14_C : bit_vector(255 downto 0) := x"7FB39A6084FEC5F9021E5AFBD7364CE2BCE97DBB5D3E443DD73A3E86DE7B047D";
   constant CPIX_NORMAL_INIT_29_BIT_00_C : bit_vector(255 downto 0) := x"C40EB3D4813860145CDF092A7C9AA7E9F9155F94B1EBDF8804EB8779C9F64B10";
   constant CPIX_NORMAL_INIT_29_BIT_01_C : bit_vector(255 downto 0) := x"131D37549C15B40EE6F06641DD8B035D99E672E7D7BF9531435826C257482605";
   constant CPIX_NORMAL_INIT_29_BIT_02_C : bit_vector(255 downto 0) := x"8A2772724949CA89C95ECABFE3B7D82B744205F63FC0D6C3618121A90135DCC8";
   constant CPIX_NORMAL_INIT_29_BIT_03_C : bit_vector(255 downto 0) := x"7C6C35ACD79CE0CAFF0FF79C3E8094429816D18C88CB840CF44AEAB7DF30185B";
   constant CPIX_NORMAL_INIT_29_BIT_04_C : bit_vector(255 downto 0) := x"1B250D6EC02029D0078FB32E59F0688575FB0479BE6827F07D268A22945E99C2";
   constant CPIX_NORMAL_INIT_29_BIT_05_C : bit_vector(255 downto 0) := x"BD54EF8AB896363C9CCBADCB0FFD52602D305A15765BA157327C9148609AE72B";
   constant CPIX_NORMAL_INIT_29_BIT_06_C : bit_vector(255 downto 0) := x"FF30B07785D5F5CCFDBDA2753A8B5AB93A4664D45C478181043059D08BEB7C97";
   constant CPIX_NORMAL_INIT_29_BIT_07_C : bit_vector(255 downto 0) := x"E787359EB9A71C571264CCE9A5449638882306532D8ECE27B397C2825B5072B1";
   constant CPIX_NORMAL_INIT_29_BIT_08_C : bit_vector(255 downto 0) := x"53D53BB753C94BF2A5466E498451E18C5458B3938C76CF36CE1EEE53246FEF77";
   constant CPIX_NORMAL_INIT_29_BIT_09_C : bit_vector(255 downto 0) := x"B8A2EE38457E0E13CBC93DA556CF07FFEA88DC3798DA5848F6DCAB3517F9CA69";
   constant CPIX_NORMAL_INIT_29_BIT_10_C : bit_vector(255 downto 0) := x"99859E239113E689F7F5C8DD86198D3394121558135A964B6A89E67F92FD1BE0";
   constant CPIX_NORMAL_INIT_29_BIT_11_C : bit_vector(255 downto 0) := x"8B8C33E0FA212DBAB7F8129BE56CF4E52C3270003CF2638056A8937FEE942EAF";
   constant CPIX_NORMAL_INIT_29_BIT_12_C : bit_vector(255 downto 0) := x"41617EFE7E6F81F42C27EB0408B4F14FF2F540E50F4492E8964C269B09FFB791";
   constant CPIX_NORMAL_INIT_29_BIT_13_C : bit_vector(255 downto 0) := x"80AED57F7EB59166CFEFB2D28DD087E08109DDFA47A2ECAE6FA5A3151981CEC5";
   constant CPIX_NORMAL_INIT_29_BIT_14_C : bit_vector(255 downto 0) := x"CF6D1AC0F3380C6F1028833C96361C8A249C443AA8F15C3AD93272D4035FFF88";
   constant CPIX_NORMAL_INIT_2A_BIT_00_C : bit_vector(255 downto 0) := x"4773AE29D8F37AC171B9FD4909AC98A30E62B4A5FEDC17663A835CE0D8B00259";
   constant CPIX_NORMAL_INIT_2A_BIT_01_C : bit_vector(255 downto 0) := x"3A202C143BD1168F7D06338CA771681B0147DE2836009F3ED20DC559BDDE87AC";
   constant CPIX_NORMAL_INIT_2A_BIT_02_C : bit_vector(255 downto 0) := x"213B4FE7E20384DD0815009948E18D4B1B16BD51B0C9CA46BF522789A9AD6888";
   constant CPIX_NORMAL_INIT_2A_BIT_03_C : bit_vector(255 downto 0) := x"92AEE600A3B6E0948866008240C4F0308DE642889C1009EDF57950E824F19A39";
   constant CPIX_NORMAL_INIT_2A_BIT_04_C : bit_vector(255 downto 0) := x"CDE7090B070F83EC5D50E5C7C900CF3DD5005CE1E386C8A8BDAE753746FBF56F";
   constant CPIX_NORMAL_INIT_2A_BIT_05_C : bit_vector(255 downto 0) := x"EE2DA6A1C37A1E5D196BDFB94E71F207E5AA95786BB7A425113326FE2CA4CD7F";
   constant CPIX_NORMAL_INIT_2A_BIT_06_C : bit_vector(255 downto 0) := x"FD5D54B99C6E17A5F38DDFFD2F337FADEA7CF39B82952E5B2B3DB9FBB41A11C7";
   constant CPIX_NORMAL_INIT_2A_BIT_07_C : bit_vector(255 downto 0) := x"9DFF418F7AF9BD8BF5BDFF35B4D9CF4D5EDB814A1341F0EBFBAE99376D423505";
   constant CPIX_NORMAL_INIT_2A_BIT_08_C : bit_vector(255 downto 0) := x"ACD44DD522B9BE76273A671FE6479D1FFFD64134AF2623179049B54BE68BBF3D";
   constant CPIX_NORMAL_INIT_2A_BIT_09_C : bit_vector(255 downto 0) := x"AE35A753D5CAFF1637CEC7D91F47B6C782635D970BA8A7F194BB873A554EA579";
   constant CPIX_NORMAL_INIT_2A_BIT_10_C : bit_vector(255 downto 0) := x"ADDB7ED441AC352A7A4C85E1FF1ECC27D9F1F337AEE913BCF30A718EE01CA315";
   constant CPIX_NORMAL_INIT_2A_BIT_11_C : bit_vector(255 downto 0) := x"9FA5CA162B72FDF6D26E87532505E09B4C96EB4928A48F219778EAA638E310B5";
   constant CPIX_NORMAL_INIT_2A_BIT_12_C : bit_vector(255 downto 0) := x"A70A5038683D96064A382759A9C77EE15A96142DB148837F45DB31B49FFC22A5";
   constant CPIX_NORMAL_INIT_2A_BIT_13_C : bit_vector(255 downto 0) := x"BBB82BC22C94D130E42E071B688F94110FBC5A645E4057D17AE3ED6EE4454809";
   constant CPIX_NORMAL_INIT_2A_BIT_14_C : bit_vector(255 downto 0) := x"2A845EC2CBD7E74E0874258B902294D358E186A8223AEA7CF8272BE09FE3E8B3";
   constant CPIX_NORMAL_INIT_2B_BIT_00_C : bit_vector(255 downto 0) := x"C16A6D7D23BD42D7F6D4B578667AB6A17989704A7BFDA6F7CD3710BE7F6C8489";
   constant CPIX_NORMAL_INIT_2B_BIT_01_C : bit_vector(255 downto 0) := x"1BA42989732D577B35A1485F5B7A18D5B7C28B20CC9E71FA3F7CD40783F78840";
   constant CPIX_NORMAL_INIT_2B_BIT_02_C : bit_vector(255 downto 0) := x"04C336B1220F9CF72114EA1DB9554CD795ADBCC19583021CFEAD0090258D0452";
   constant CPIX_NORMAL_INIT_2B_BIT_03_C : bit_vector(255 downto 0) := x"F61BAADC1CE81FDC3B58D49A0C6E872A92C42425BCBD0F735B5E0B4A804BF44F";
   constant CPIX_NORMAL_INIT_2B_BIT_04_C : bit_vector(255 downto 0) := x"5F0453CD37C64FBDEA009BC7E88C1293A2F60141E2C45757B88C8E97E51AF044";
   constant CPIX_NORMAL_INIT_2B_BIT_05_C : bit_vector(255 downto 0) := x"F196F716C02ABF4FD298C57216D24ECF796C2C0BA575509E2A2555BE7DA91EA5";
   constant CPIX_NORMAL_INIT_2B_BIT_06_C : bit_vector(255 downto 0) := x"D915392D87DB5FEB2B872588F0D934AF5E29159EA9F0955264CDC19DB294028D";
   constant CPIX_NORMAL_INIT_2B_BIT_07_C : bit_vector(255 downto 0) := x"52231F2D379D51BDAF480867B2E6B7D165D7B2169F71B627129B3B893A0CB5FF";
   constant CPIX_NORMAL_INIT_2B_BIT_08_C : bit_vector(255 downto 0) := x"7CF6B3021BC3EF2C8380730D3FEDA9056098C03A32FF94EFBA779F7427790734";
   constant CPIX_NORMAL_INIT_2B_BIT_09_C : bit_vector(255 downto 0) := x"BC10BF9AAE99C181B6BE8F5185E10C9FD32563CF19A83A54D93B9FF120058FF0";
   constant CPIX_NORMAL_INIT_2B_BIT_10_C : bit_vector(255 downto 0) := x"B6D6B9A9190F129D2D13737CB9AD23CE0DC04E2530B2392084FD030FACD29C92";
   constant CPIX_NORMAL_INIT_2B_BIT_11_C : bit_vector(255 downto 0) := x"B80B5D51F214CB65FBCAF0F66A41C7DAACB6D47B831F2CD2799BBF05151D81B8";
   constant CPIX_NORMAL_INIT_2B_BIT_12_C : bit_vector(255 downto 0) := x"9058EBF96E8AD4F0AD27A8C000BF3C6C6DBCD246E69973CB9847CD3A660A45F2";
   constant CPIX_NORMAL_INIT_2B_BIT_13_C : bit_vector(255 downto 0) := x"1E75DA5530377CCE82BCB25D178C60B4AAFC3FE07C8567069D03E8AF8631A02A";
   constant CPIX_NORMAL_INIT_2B_BIT_14_C : bit_vector(255 downto 0) := x"043056DA14E44BC0A587113A1D20EC18974252D3BF41CF153FB6C57DA5E2D91C";
   constant CPIX_NORMAL_INIT_2C_BIT_00_C : bit_vector(255 downto 0) := x"D9EE592D6C138137CA8F664E703D19F82D57DF376DDA1164924607E6D46050EB";
   constant CPIX_NORMAL_INIT_2C_BIT_01_C : bit_vector(255 downto 0) := x"3B66C0C454E028DF809E5CDFB33B5A4A2FFB51A884C47A0065DBED9F341391B3";
   constant CPIX_NORMAL_INIT_2C_BIT_02_C : bit_vector(255 downto 0) := x"57EE826BDFE5A829BB2F2360340DA1F95AB8671EE39F96F2B408BDA0E6C98816";
   constant CPIX_NORMAL_INIT_2C_BIT_03_C : bit_vector(255 downto 0) := x"2FD0A3C1A97780528C8A18FB83A6B03EFE8E860FF7CAF19479F96B6682E83335";
   constant CPIX_NORMAL_INIT_2C_BIT_04_C : bit_vector(255 downto 0) := x"52722CBEF28C66C6D46C97DE98E783FFD134C3E7E2E5DAB33D99EE28CA2EA902";
   constant CPIX_NORMAL_INIT_2C_BIT_05_C : bit_vector(255 downto 0) := x"081182948278D6E1076303011A9571126F7D9BE17E10DAA7A6E355FC9DB4E7EF";
   constant CPIX_NORMAL_INIT_2C_BIT_06_C : bit_vector(255 downto 0) := x"AF7475423B063A47D126CC499C49DF63D6D7C250302DE122A6868A98D648730D";
   constant CPIX_NORMAL_INIT_2C_BIT_07_C : bit_vector(255 downto 0) := x"264B6690F68B59B780DBB275928430C7C49D12B8402095643A95216B753931BF";
   constant CPIX_NORMAL_INIT_2C_BIT_08_C : bit_vector(255 downto 0) := x"D8D19272C373295D9A41B9B9091B254ECE960171C1B73201CCAEE5FB2A79E96A";
   constant CPIX_NORMAL_INIT_2C_BIT_09_C : bit_vector(255 downto 0) := x"B76B9CC504337451FC011353DB7BC60B02FE62AC60C4830F1A22F3BFDDFB24A6";
   constant CPIX_NORMAL_INIT_2C_BIT_10_C : bit_vector(255 downto 0) := x"76E06D48D7179B6FE66E2E5D22427B3BFCF097E2DB6D2838BC435BC0D48F0858";
   constant CPIX_NORMAL_INIT_2C_BIT_11_C : bit_vector(255 downto 0) := x"89B7D601F8CF149970B79BD184E267A5A6296D41040755E1D24826A9763336E4";
   constant CPIX_NORMAL_INIT_2C_BIT_12_C : bit_vector(255 downto 0) := x"366DB662E3C6AD933DA0D7A344D7909CC35621B000A0D4522B64C7415F59009A";
   constant CPIX_NORMAL_INIT_2C_BIT_13_C : bit_vector(255 downto 0) := x"9C43B1CFC42822DF7F5258E63CD0D5D392A4453E60158425D8B602EEE43494D0";
   constant CPIX_NORMAL_INIT_2C_BIT_14_C : bit_vector(255 downto 0) := x"2CB1F995FADDA5FCD70E03AF69353D2F3892EF0FFFDE28FC354F7CEBAC8BDBC4";
   constant CPIX_NORMAL_INIT_2D_BIT_00_C : bit_vector(255 downto 0) := x"0BBDB263100CD06561172A6AED0034582F55BE1139F337811656235817776155";
   constant CPIX_NORMAL_INIT_2D_BIT_01_C : bit_vector(255 downto 0) := x"83427640083D130105918DC6BF0D33BDE61F8AF30B16EE67DA445DF04E882F83";
   constant CPIX_NORMAL_INIT_2D_BIT_02_C : bit_vector(255 downto 0) := x"A4B4E6FE871CB399C4BD4F137BD466690F2DFAE78229F18D6319E09D39BAA3DC";
   constant CPIX_NORMAL_INIT_2D_BIT_03_C : bit_vector(255 downto 0) := x"4EC8A79B6B0E058434BEFF882A16ED018C7DBAE8427F59B36CCE17538D5A30F9";
   constant CPIX_NORMAL_INIT_2D_BIT_04_C : bit_vector(255 downto 0) := x"C4116CF80B1D85B6C62A4C250DE262A72B50CB18E548E122474189990304EB9F";
   constant CPIX_NORMAL_INIT_2D_BIT_05_C : bit_vector(255 downto 0) := x"5F51F80D5578D782A290B90C64E838F34AFC2387D75F0D21E3E1C2825CE4D91C";
   constant CPIX_NORMAL_INIT_2D_BIT_06_C : bit_vector(255 downto 0) := x"2D4BBF54C03EDECFA48BC163DAA3355CA2B4D4419B79E86E90CF27058162E058";
   constant CPIX_NORMAL_INIT_2D_BIT_07_C : bit_vector(255 downto 0) := x"CF7403C139C3E7F9B231E814EC6547344C653F75EDBBC48F1E7FE5766AD7A535";
   constant CPIX_NORMAL_INIT_2D_BIT_08_C : bit_vector(255 downto 0) := x"4D5424C6706B38C451EC8266EA5530B2B237E65077F5951D922967E6DBFA575B";
   constant CPIX_NORMAL_INIT_2D_BIT_09_C : bit_vector(255 downto 0) := x"D1C742F3481A210F4D5C2C31DBE6375F4263588F1C583A4A06DB74B80BEF8700";
   constant CPIX_NORMAL_INIT_2D_BIT_10_C : bit_vector(255 downto 0) := x"ACA4F52D5DC2088827A637F00E9E6B6B68F982607A9F22FA6A3BF885AE3EE2CA";
   constant CPIX_NORMAL_INIT_2D_BIT_11_C : bit_vector(255 downto 0) := x"18763FE87E9D01FAF9C14B2EC575B4DBD262221162C313B1C6BA354CFFC388F8";
   constant CPIX_NORMAL_INIT_2D_BIT_12_C : bit_vector(255 downto 0) := x"09FE7F01BA59D76637C986F8A1ACC5D07DD04310184FF829A3396A3DBD02165D";
   constant CPIX_NORMAL_INIT_2D_BIT_13_C : bit_vector(255 downto 0) := x"5E5892B2317DD50E0453B5DD7D7C20EE09DF7DEEF60AC70FE3DC6151A66667FE";
   constant CPIX_NORMAL_INIT_2D_BIT_14_C : bit_vector(255 downto 0) := x"9669E7996BE0AA526F29E2341963E8D5BC7D3DFD0744620739E07F1986CFCB8D";
   constant CPIX_NORMAL_INIT_2E_BIT_00_C : bit_vector(255 downto 0) := x"57D5455E9521E9EAFED7AB47AD13F648C3B64B16C375D8F0FADF8FFE50502809";
   constant CPIX_NORMAL_INIT_2E_BIT_01_C : bit_vector(255 downto 0) := x"99E6BA9AE78B71FEB4D30FB33C52E2A2B2B2ED6C50ACAB6979B4651F2A9A5C7A";
   constant CPIX_NORMAL_INIT_2E_BIT_02_C : bit_vector(255 downto 0) := x"0A218BAE7211C7CD147A2E7A01A008F25F5EE0F26212315DA903E52C28068C56";
   constant CPIX_NORMAL_INIT_2E_BIT_03_C : bit_vector(255 downto 0) := x"66CD90388DE3DE06B6E39D20BCE8E5BB440B07C90C9D1378D0C01DF93F3BB9B1";
   constant CPIX_NORMAL_INIT_2E_BIT_04_C : bit_vector(255 downto 0) := x"F9CA5473604C42665FEF349FD1CF153BF7BA82CE1DC4FB4666458CB074412657";
   constant CPIX_NORMAL_INIT_2E_BIT_05_C : bit_vector(255 downto 0) := x"7D75CC34D849B80C77AACD6F01BFC0BA02C1D3F49BA3E8744D00F1BA794E7979";
   constant CPIX_NORMAL_INIT_2E_BIT_06_C : bit_vector(255 downto 0) := x"CE1C3A753AA8E353AA5EA78DD04850C05FB14460DD27BC4F8E9F032296DCFBB1";
   constant CPIX_NORMAL_INIT_2E_BIT_07_C : bit_vector(255 downto 0) := x"723CB73169EEB8C4A884528681308F15FA3F003897D6691CB2356F5BDF67E607";
   constant CPIX_NORMAL_INIT_2E_BIT_08_C : bit_vector(255 downto 0) := x"D8CA2E393A468CE2299D2895C048538FC21977739B9CD32DD890308DA6C267C5";
   constant CPIX_NORMAL_INIT_2E_BIT_09_C : bit_vector(255 downto 0) := x"7253E3D2149F797C5E6837758B650CE9B6ECA7E35930CA492E84F1ACB8ABF115";
   constant CPIX_NORMAL_INIT_2E_BIT_10_C : bit_vector(255 downto 0) := x"C834FF8D480108DD8F79403545F735E61CF35805BE907DE166FAE8F3BF8ABF5C";
   constant CPIX_NORMAL_INIT_2E_BIT_11_C : bit_vector(255 downto 0) := x"1FF3FA313B0C72541FD3E846779D65D2C3367A10EB2E26C9F12267DF1D0D10D8";
   constant CPIX_NORMAL_INIT_2E_BIT_12_C : bit_vector(255 downto 0) := x"727253AFE6D8CD3736D2F6EA95AE24EEC260C028B0BF37D308FF37A081BAF5A2";
   constant CPIX_NORMAL_INIT_2E_BIT_13_C : bit_vector(255 downto 0) := x"D88080947AD5FF24165D82D08B65FFED48EBC9FFBCC2336CC33C0204327BA12E";
   constant CPIX_NORMAL_INIT_2E_BIT_14_C : bit_vector(255 downto 0) := x"723E830B9A6027D58ECB8E8D24F93C76E2691F2FEA94286E71BA95C804875AA4";
   constant CPIX_NORMAL_INIT_2F_BIT_00_C : bit_vector(255 downto 0) := x"59A0E4E56570FC742F3C5F09ED5F9BE5625A6ED9DAF9FB4B894A08921B498351";
   constant CPIX_NORMAL_INIT_2F_BIT_01_C : bit_vector(255 downto 0) := x"17D4AF2C47839697798B2312C19787785ECE1FAC17254430DE9CD40834C4A1AC";
   constant CPIX_NORMAL_INIT_2F_BIT_02_C : bit_vector(255 downto 0) := x"A0C111B5AD16873DAA6991110EF31C6E29E7ACE9289E041CB7067C17DEE23DC0";
   constant CPIX_NORMAL_INIT_2F_BIT_03_C : bit_vector(255 downto 0) := x"F97BA5DCF00DB29B7244FC9EC18FF701AC533910179E01A34C00BA5518F271BF";
   constant CPIX_NORMAL_INIT_2F_BIT_04_C : bit_vector(255 downto 0) := x"C3E3DBF30A80E3CA6799A0374D68D5E1423FA5DBDBE4B3D6C9A7F21D999ED127";
   constant CPIX_NORMAL_INIT_2F_BIT_05_C : bit_vector(255 downto 0) := x"D9936AA91E870DBC15F94BB31449EDD2B7E4CA02E43A16DA123FFC5DCD0FD193";
   constant CPIX_NORMAL_INIT_2F_BIT_06_C : bit_vector(255 downto 0) := x"93ADF88D000D67E14CBB90E72E7EB12B34AC8D37372FBED907613CB7F3BC3AF9";
   constant CPIX_NORMAL_INIT_2F_BIT_07_C : bit_vector(255 downto 0) := x"85C9E8B2CC34A6FD0647F7F100F4F509CCD78D9F9825D1CDCB850D29567F9B09";
   constant CPIX_NORMAL_INIT_2F_BIT_08_C : bit_vector(255 downto 0) := x"051FFF0C97D3613A7ED9249506042816E2031A39350CAE5399F6DF15A2D49F28";
   constant CPIX_NORMAL_INIT_2F_BIT_09_C : bit_vector(255 downto 0) := x"16D913AACC0164AED2511513FE8354F07E94FBD292055EA9978C484F1CC0AAE9";
   constant CPIX_NORMAL_INIT_2F_BIT_10_C : bit_vector(255 downto 0) := x"3AB12F3A93A9C974B071144D52F63823CEADB2450E20D7B3AC8F6CF01A4B1F01";
   constant CPIX_NORMAL_INIT_2F_BIT_11_C : bit_vector(255 downto 0) := x"329556CC0ECA5A1D854FB3CB6F8926A533B9841A22A9C7AA9188367D4118A369";
   constant CPIX_NORMAL_INIT_2F_BIT_12_C : bit_vector(255 downto 0) := x"34698E0A2F2F9606B75E18575D57700F81969F3498685AFCB563A94A33D584E4";
   constant CPIX_NORMAL_INIT_2F_BIT_13_C : bit_vector(255 downto 0) := x"2485171229FBA7017D0D94302B2327A92AB928EC2697A3B90B9175A0536C9FFE";
   constant CPIX_NORMAL_INIT_2F_BIT_14_C : bit_vector(255 downto 0) := x"06E481A42CB14E608FC781B6B9EDBC34CA65612C5DD6CB86C30C98717D246CA0";
   constant CPIX_NORMAL_INIT_30_BIT_00_C : bit_vector(255 downto 0) := x"54670A94896083502022AF7D553C41BA39430B08CF5AE86E85C1C6461D3436BD";
   constant CPIX_NORMAL_INIT_30_BIT_01_C : bit_vector(255 downto 0) := x"968F1A5620DA4B0424E5C696233646025BE2769979F4978E8F3A1B9847E4B1CC";
   constant CPIX_NORMAL_INIT_30_BIT_02_C : bit_vector(255 downto 0) := x"39454C0F77C56271AF410E004E737FDBF9E58A76958BDE1E20273CCDDE7663A3";
   constant CPIX_NORMAL_INIT_30_BIT_03_C : bit_vector(255 downto 0) := x"C9433DC951792465D1E2637E9B56A13C521A251E17725A09981BE011E83E63F3";
   constant CPIX_NORMAL_INIT_30_BIT_04_C : bit_vector(255 downto 0) := x"0A05F34F5285A08B37AEA155C6F8F2A075469038C09C359E5C9E5E07EE6B401A";
   constant CPIX_NORMAL_INIT_30_BIT_05_C : bit_vector(255 downto 0) := x"F04C2BFC7DD41C5F87F553C7F3B95904184397617CBFEFE83FFAA9BDF3329139";
   constant CPIX_NORMAL_INIT_30_BIT_06_C : bit_vector(255 downto 0) := x"9AE2C51AD006699418E0F2DA7E83D06E592BC35EAB6A7A648B796CD9EACED96F";
   constant CPIX_NORMAL_INIT_30_BIT_07_C : bit_vector(255 downto 0) := x"CA6F58D872298D014A1CCCAF6D1052778F3B29638E3F102504F7E8C178FFD7B1";
   constant CPIX_NORMAL_INIT_30_BIT_08_C : bit_vector(255 downto 0) := x"957C158ED0365B309332E98D7B77B635C474561A4B57BAC3D338560D4752F838";
   constant CPIX_NORMAL_INIT_30_BIT_09_C : bit_vector(255 downto 0) := x"C685FA3268F86ADE5953EA73F2B575DFDB87912711F59C1F823A832ED05A25BE";
   constant CPIX_NORMAL_INIT_30_BIT_10_C : bit_vector(255 downto 0) := x"9A3F1B20EFCA8AFDC7E17A1F13EA88EA99A7A74C142ED33942AA54C661C37666";
   constant CPIX_NORMAL_INIT_30_BIT_11_C : bit_vector(255 downto 0) := x"3767CA16AB88DCAEE4BC033AFCBCD2456319A574A2F54A132CB7493C55348926";
   constant CPIX_NORMAL_INIT_30_BIT_12_C : bit_vector(255 downto 0) := x"C676BE9D2DD8C58E1F4EE5514FAE80C52F4F9BD36BC974EB6EA2CCAA3C0F14FA";
   constant CPIX_NORMAL_INIT_30_BIT_13_C : bit_vector(255 downto 0) := x"9101F8A638FF03BEAA046CF655D6BFF053D0632CA8DFE124F84B6164772D2628";
   constant CPIX_NORMAL_INIT_30_BIT_14_C : bit_vector(255 downto 0) := x"CE356BC743CA19BDE79B9928DBD03CF59850BD8AF84812153D415AF353CC29CC";
   constant CPIX_NORMAL_INIT_31_BIT_00_C : bit_vector(255 downto 0) := x"C41877ED0F65ABDFF16B151188D1AD538190D7677F0DD2786263CC8D299E472C";
   constant CPIX_NORMAL_INIT_31_BIT_01_C : bit_vector(255 downto 0) := x"1F69A86288EC6908965E9FF249C34591093DF811C691D23F9226A70557D13115";
   constant CPIX_NORMAL_INIT_31_BIT_02_C : bit_vector(255 downto 0) := x"6B5B630D8BEEA259EAB10B5E361FCF50E55E07BDC1635C9B715C734839518C1C";
   constant CPIX_NORMAL_INIT_31_BIT_03_C : bit_vector(255 downto 0) := x"91B929042E39E57ADDAE23998E4241D5CF3DEB9F0166DDF219724E77FEA1614E";
   constant CPIX_NORMAL_INIT_31_BIT_04_C : bit_vector(255 downto 0) := x"7D23D0DB9A9B77A25FCE40FB1F9E5D53451A681A63FE0FC573E0D01C3673A0B9";
   constant CPIX_NORMAL_INIT_31_BIT_05_C : bit_vector(255 downto 0) := x"CF1075114B791FA7BECBBA31B1F62087BFFDF5145803A4285744363A349CAB19";
   constant CPIX_NORMAL_INIT_31_BIT_06_C : bit_vector(255 downto 0) := x"398FCD509F83A39B13E6C2F0234780468A9D8462C034170DFFF9A4A348B644D4";
   constant CPIX_NORMAL_INIT_31_BIT_07_C : bit_vector(255 downto 0) := x"B3A4A3A2D24DD9E50C0B6A94F63F7AEA8B4E2840A272602654A74D07C572C3AC";
   constant CPIX_NORMAL_INIT_31_BIT_08_C : bit_vector(255 downto 0) := x"BB8859F2D8430D5200CEA6C7EB3DC2659FE8406152D1E75940736C30A6A006A3";
   constant CPIX_NORMAL_INIT_31_BIT_09_C : bit_vector(255 downto 0) := x"ACE46C10BDBF5398075820F412929DE40F5C2C80B748EF4690A684F706AA19FF";
   constant CPIX_NORMAL_INIT_31_BIT_10_C : bit_vector(255 downto 0) := x"597B118A1FF5624CD623C55DDFD400F0D3C752F78D90B1ABCCBCF684AEF7F0CE";
   constant CPIX_NORMAL_INIT_31_BIT_11_C : bit_vector(255 downto 0) := x"1EDE273EAABABCA3879A13AFC56642C740A8A128C6CE4197CFA7E9C9DD3A8061";
   constant CPIX_NORMAL_INIT_31_BIT_12_C : bit_vector(255 downto 0) := x"3F2EACB7698903BE62740A0B1C73A28AAE408640B210A0C4716F0BA8ED2944FE";
   constant CPIX_NORMAL_INIT_31_BIT_13_C : bit_vector(255 downto 0) := x"9247ACF2FAD06BA8EBA0EFCDC43DFDB009580820CA8B0D43F6C2A78A80B46DAB";
   constant CPIX_NORMAL_INIT_31_BIT_14_C : bit_vector(255 downto 0) := x"003D56C434A1CA7C713EB9BD28247BFB573D5B9F5587D5BAAC747C60DBD9FB68";
   constant CPIX_NORMAL_INIT_32_BIT_00_C : bit_vector(255 downto 0) := x"F92030B4D422D357E73EEBD6252EF79C05F14E0C40FBDD0760AF9EE5DDFF94E6";
   constant CPIX_NORMAL_INIT_32_BIT_01_C : bit_vector(255 downto 0) := x"417195F92154A2C1BA5A825108F08E62C7E8938C1F28676C5CFC4B21381B012F";
   constant CPIX_NORMAL_INIT_32_BIT_02_C : bit_vector(255 downto 0) := x"A43D30BB361D026BAF773DFD38B9F5B1FCCEA5FD8A9F61B03D75B47FB235AC75";
   constant CPIX_NORMAL_INIT_32_BIT_03_C : bit_vector(255 downto 0) := x"242E5FAC3EEC25648C079462F8BFFC931E1308B392B2DF9B7E1F040EAB912BDA";
   constant CPIX_NORMAL_INIT_32_BIT_04_C : bit_vector(255 downto 0) := x"E385492C691CCB969C87853FDE459DF618079C20D17CEBB552A8263D7F7F8399";
   constant CPIX_NORMAL_INIT_32_BIT_05_C : bit_vector(255 downto 0) := x"7CACCF5D039638DFA8A8EADF0B882C2B6A21F29E1601CB634711A6C120217612";
   constant CPIX_NORMAL_INIT_32_BIT_06_C : bit_vector(255 downto 0) := x"BFEB60ED26B68930D9A0778CC50AF4015489B1AA252A7869B9E5B5370BBA4C5F";
   constant CPIX_NORMAL_INIT_32_BIT_07_C : bit_vector(255 downto 0) := x"5626E2C29BE914775E31AC1C2D912D0914AD0C18B266CD0608F926887D8A6F3D";
   constant CPIX_NORMAL_INIT_32_BIT_08_C : bit_vector(255 downto 0) := x"104950502DAE646F9A7F38615033FECF8226BEC94CED9E1D6CBCCDA9A1C47FB6";
   constant CPIX_NORMAL_INIT_32_BIT_09_C : bit_vector(255 downto 0) := x"51111FE64686A2CF02AD80BDE547A839D16B909323F5729FB16A2BBEAE2CD253";
   constant CPIX_NORMAL_INIT_32_BIT_10_C : bit_vector(255 downto 0) := x"FBB48F9CCDDA99F0467835F049071D07069A04960BC6CE34EBB1363D263D1433";
   constant CPIX_NORMAL_INIT_32_BIT_11_C : bit_vector(255 downto 0) := x"01B5C0A8D6998B9714C1B83F7BAD80255602E1CADB7C2E5E6336C9D9D0586105";
   constant CPIX_NORMAL_INIT_32_BIT_12_C : bit_vector(255 downto 0) := x"A079D7EF961CCC685B856957FAD26EF3CBE0018C3F2F479F5C05EC40DCC1DFE0";
   constant CPIX_NORMAL_INIT_32_BIT_13_C : bit_vector(255 downto 0) := x"27D713DB634324DEA9C798CCF9786DD620DBDD4C31AD6A6CBD872189DBC3AE51";
   constant CPIX_NORMAL_INIT_32_BIT_14_C : bit_vector(255 downto 0) := x"F7C7A3D9AEC89714A60E0AFFBE78F7FB4B5896E12E1FCB430055154FE2F811FD";
   constant CPIX_NORMAL_INIT_33_BIT_00_C : bit_vector(255 downto 0) := x"5B07708B39909D7041ADFE2104123BCDEB94D3606C4B6ED91C44EAAF6859AF13";
   constant CPIX_NORMAL_INIT_33_BIT_01_C : bit_vector(255 downto 0) := x"9DC8290270CDFCE5C479113B643FF4BD38341291ECE933111FADC3BDE4980AAA";
   constant CPIX_NORMAL_INIT_33_BIT_02_C : bit_vector(255 downto 0) := x"255E9940FC8AD80AE30206FCBED451793AE0B0BD6A04E1A9FA2220A0D79FED34";
   constant CPIX_NORMAL_INIT_33_BIT_03_C : bit_vector(255 downto 0) := x"C6B53DEE1E7D8596A694CCB15AEC4885391F3509526781FD1C10D6C06F21D017";
   constant CPIX_NORMAL_INIT_33_BIT_04_C : bit_vector(255 downto 0) := x"4749466126D9C0FABED237E63751DF385B1566F8791411A64D5645FED32ACB56";
   constant CPIX_NORMAL_INIT_33_BIT_05_C : bit_vector(255 downto 0) := x"A8463830216566EDFE882E9C5C438BEABECE2E9C21FD5EC67929891275948A6B";
   constant CPIX_NORMAL_INIT_33_BIT_06_C : bit_vector(255 downto 0) := x"BA32B59DE33B21CC6FB12F8367CAA456C03370BD66A667F0A0FFF87E4D6E09B9";
   constant CPIX_NORMAL_INIT_33_BIT_07_C : bit_vector(255 downto 0) := x"847EAB3E6DAE1C5521B64996362FCEA89791E53ED42E3ED7EB6FB8A9923BA5FB";
   constant CPIX_NORMAL_INIT_33_BIT_08_C : bit_vector(255 downto 0) := x"DF07F8A65921E8457E4F2A7C4BFB0610FF404E55C57B6433663C3EAD43CFBB89";
   constant CPIX_NORMAL_INIT_33_BIT_09_C : bit_vector(255 downto 0) := x"521FA13D2138321F96EF33203186ED67042A6344ACF9267B6DBD4DAEA50F666D";
   constant CPIX_NORMAL_INIT_33_BIT_10_C : bit_vector(255 downto 0) := x"4F730B327994EA280B34178947429888B3672BFDCA25ED17D8E99C1FA95ADBB9";
   constant CPIX_NORMAL_INIT_33_BIT_11_C : bit_vector(255 downto 0) := x"54AAB807D09DCF97F72F233A2E8886499FB530405562DDDF8CADC72876CB9E6F";
   constant CPIX_NORMAL_INIT_33_BIT_12_C : bit_vector(255 downto 0) := x"02F5831C0FDA51691C59A71CC3B68C589F7A2E933B646BB892BCD1A1DA0F821D";
   constant CPIX_NORMAL_INIT_33_BIT_13_C : bit_vector(255 downto 0) := x"1AA7DD6229404A553471446DD90C71D53BC6A38EC830FCE6CC3C02305B437557";
   constant CPIX_NORMAL_INIT_33_BIT_14_C : bit_vector(255 downto 0) := x"029EB1CA301926297FF9BAC9702D878F915DDA54356171631A380743BF9D9504";
   constant CPIX_NORMAL_INIT_34_BIT_00_C : bit_vector(255 downto 0) := x"E8CD4FF6856B6F12443A4879856D908E666789B96113CBBF09F86A41494F45E7";
   constant CPIX_NORMAL_INIT_34_BIT_01_C : bit_vector(255 downto 0) := x"AED0890D5E73BEB332DA8E9EE2AED3793E57C087CD5DA33DBD4108022FDDBFA2";
   constant CPIX_NORMAL_INIT_34_BIT_02_C : bit_vector(255 downto 0) := x"DCD77A8DA743D3AB3E37D92DAD329B49471561FD261F22343E0E33EC87279D59";
   constant CPIX_NORMAL_INIT_34_BIT_03_C : bit_vector(255 downto 0) := x"0C107F745524D9DC47018793D7CEC41D12C261E57587E8B0AA014AF7E9139E07";
   constant CPIX_NORMAL_INIT_34_BIT_04_C : bit_vector(255 downto 0) := x"EE62491B6FCAC86912441C871E8490CB4CC25499020E134CF12EDC3B4665B97D";
   constant CPIX_NORMAL_INIT_34_BIT_05_C : bit_vector(255 downto 0) := x"705C0273F354806BB520CE30DEAB44306B45592479788386FDD9D0EB70AD7B4A";
   constant CPIX_NORMAL_INIT_34_BIT_06_C : bit_vector(255 downto 0) := x"974D0E6057247FD762D8897762E227AB7C8A606323F084B2B598C2844B41560E";
   constant CPIX_NORMAL_INIT_34_BIT_07_C : bit_vector(255 downto 0) := x"2EC15F52E3B5F3731BB841A3CB338154ED50507251496DF55898E5A10CB7C323";
   constant CPIX_NORMAL_INIT_34_BIT_08_C : bit_vector(255 downto 0) := x"90052E3026707C8F899EA73DF19C6D507F2356D313B97A7C67C14995EB29BA33";
   constant CPIX_NORMAL_INIT_34_BIT_09_C : bit_vector(255 downto 0) := x"8A022DD2F5EF5CD149DD0DE61C7F7E44A2C4147155323F737824C511C26EE26E";
   constant CPIX_NORMAL_INIT_34_BIT_10_C : bit_vector(255 downto 0) := x"C532B6760EBF5E1F55FDB4AC9C46CFAF5C1C7BDA82DFDDBA1192A4785D229CF2";
   constant CPIX_NORMAL_INIT_34_BIT_11_C : bit_vector(255 downto 0) := x"DF64493A18DB30F0823F292D694CB1EA9BB9FFFFDD0ECE3D70AAFAEE973B1C2A";
   constant CPIX_NORMAL_INIT_34_BIT_12_C : bit_vector(255 downto 0) := x"FADC247DEEBBD645C73CD49CA23DD5AD9C39FB8D6C66C23AE66FCB984D43D989";
   constant CPIX_NORMAL_INIT_34_BIT_13_C : bit_vector(255 downto 0) := x"77B0C8FF93EF192EE3308429C58F824F3C3EEBBC09F28B9C0758873BBDF739D4";
   constant CPIX_NORMAL_INIT_34_BIT_14_C : bit_vector(255 downto 0) := x"009D7EA177FA022821531F5F0E05BE2F1CCC6BBA37EAFD1F5D8290999E20FBA1";
   constant CPIX_NORMAL_INIT_35_BIT_00_C : bit_vector(255 downto 0) := x"C412DFFF0725AB8FBAB51D32A68B0687CA15F8215FDB40DF2E358D5B5020A2A5";
   constant CPIX_NORMAL_INIT_35_BIT_01_C : bit_vector(255 downto 0) := x"C0EBDEEDB172600261F725A7000475C0737B8B2A93FCD44FAE632C8F1C4954E6";
   constant CPIX_NORMAL_INIT_35_BIT_02_C : bit_vector(255 downto 0) := x"DBF0B805A4D72AB80711ECA66AC3416E5C2812E5ECBDB57BEE2317D9D574D832";
   constant CPIX_NORMAL_INIT_35_BIT_03_C : bit_vector(255 downto 0) := x"F48614946FFD86A0A4F7E84EA606B857C3066C62A9F95DD352D95641FA3BC7F2";
   constant CPIX_NORMAL_INIT_35_BIT_04_C : bit_vector(255 downto 0) := x"C01A755101A39F6BA7A8208315F754E29F144759450AB0A872D0AE8DA6D06A97";
   constant CPIX_NORMAL_INIT_35_BIT_05_C : bit_vector(255 downto 0) := x"CF8ADA7CF1B513849A187E0F1286C9FD732B6D7BE321B73FE5AC9D43E0968227";
   constant CPIX_NORMAL_INIT_35_BIT_06_C : bit_vector(255 downto 0) := x"969CEEB4D071ADCCB7834172E568C4895A63B2D5EF7B56499FD0788265387794";
   constant CPIX_NORMAL_INIT_35_BIT_07_C : bit_vector(255 downto 0) := x"0FE6F56C65524D6FC21FFBF5A915C3493D96DB07D2FB905BF76E2F401A26D511";
   constant CPIX_NORMAL_INIT_35_BIT_08_C : bit_vector(255 downto 0) := x"F8BD0E762651251BF1546F320103C4E0C31D077BF3BFCD2B50E98FEFA2EFB1A9";
   constant CPIX_NORMAL_INIT_35_BIT_09_C : bit_vector(255 downto 0) := x"8B2AC6D80DB6E0D141E718A6BA82551BA8EB5126EBEF32AE2E3F30D883C8B0FA";
   constant CPIX_NORMAL_INIT_35_BIT_10_C : bit_vector(255 downto 0) := x"2134DAE2719F9A8BF8EC041CADF0A48CC595B0DAB66F191562DAA2345D571C34";
   constant CPIX_NORMAL_INIT_35_BIT_11_C : bit_vector(255 downto 0) := x"79CB2230859E463C6C1E00B8664BAE2B2512E63CD36CC691428F889F1C3B4E0D";
   constant CPIX_NORMAL_INIT_35_BIT_12_C : bit_vector(255 downto 0) := x"AFDD71871BAF066263A6841BE6AD42680AC7D86A8726719D3DD55CE62CD25443";
   constant CPIX_NORMAL_INIT_35_BIT_13_C : bit_vector(255 downto 0) := x"E2E21C2717C7195187BD7B4F999A775ED75D6F980CE6DA3C7DCA2BD38C801F5D";
   constant CPIX_NORMAL_INIT_35_BIT_14_C : bit_vector(255 downto 0) := x"DAD75D4E43BB352DA091FD2D97D73DE9ACCA8BF967622148C31EE2168E4EAFBB";
   constant CPIX_NORMAL_INIT_36_BIT_00_C : bit_vector(255 downto 0) := x"63322C65C88505B54294B61E85723EF8BD96B52DE6204C8042DDC3C82FC3F640";
   constant CPIX_NORMAL_INIT_36_BIT_01_C : bit_vector(255 downto 0) := x"1F1B7054AD9837788D1D4E5AE0B91C89C5E6020A3DDD28BE39C0754E01CA2E32";
   constant CPIX_NORMAL_INIT_36_BIT_02_C : bit_vector(255 downto 0) := x"1BC4C2A1A8D4B34ED32C60F23D23E32735CAA320330F98496FC3058D5361A50E";
   constant CPIX_NORMAL_INIT_36_BIT_03_C : bit_vector(255 downto 0) := x"4EB9C6CA08125B5B3DD10270988C3E32CA27C689CCEB8AF87108D3B520549C06";
   constant CPIX_NORMAL_INIT_36_BIT_04_C : bit_vector(255 downto 0) := x"BD4C8436F6573C30238EE869887C874DA8B8E7F155F66D34E3CE869C549843FA";
   constant CPIX_NORMAL_INIT_36_BIT_05_C : bit_vector(255 downto 0) := x"5658219E90C9A84A943523A544AA538447B8750CF51210A2C285F2685FD12E92";
   constant CPIX_NORMAL_INIT_36_BIT_06_C : bit_vector(255 downto 0) := x"58D045E630083879F38A1A8BEF12809331AB1E5C9C3A8873284567A725091127";
   constant CPIX_NORMAL_INIT_36_BIT_07_C : bit_vector(255 downto 0) := x"5A71EA380059E2C3FB54D0E6A401832CDF5EBF42C3BAE72B459C41F942798DC4";
   constant CPIX_NORMAL_INIT_36_BIT_08_C : bit_vector(255 downto 0) := x"E98FAE257D341B4E7A6266346B76A190D1D2BAF40F436FE70275822AF417E438";
   constant CPIX_NORMAL_INIT_36_BIT_09_C : bit_vector(255 downto 0) := x"6344716B4FAD5F862C5215C02E7F6A6551C79AFF3D5C051CEC93EB79C1075713";
   constant CPIX_NORMAL_INIT_36_BIT_10_C : bit_vector(255 downto 0) := x"E2D2051F3EBEA7D2447BCD1FBFFFC62A8468573078A7B73E0DBC58FD49907C33";
   constant CPIX_NORMAL_INIT_36_BIT_11_C : bit_vector(255 downto 0) := x"BD999CCFBFA686670FCAB65BC0543F1A97CACBEB49958741F29D0DC8D3CD34DD";
   constant CPIX_NORMAL_INIT_36_BIT_12_C : bit_vector(255 downto 0) := x"805961951DE67A05D66C4DFA7BF79CC858B6A4453E521FEAF148A14BFBEDC2AE";
   constant CPIX_NORMAL_INIT_36_BIT_13_C : bit_vector(255 downto 0) := x"6EE229C28DAD425F3CD3ED8B952DD1AD61B553C3C35335C2603E02A6157E151E";
   constant CPIX_NORMAL_INIT_36_BIT_14_C : bit_vector(255 downto 0) := x"25F29739AC545261733E885E683FCB884287582FCBDA2C717954DEE0D1832185";
   constant CPIX_NORMAL_INIT_37_BIT_00_C : bit_vector(255 downto 0) := x"4E6A50FF1EB7F1495CFFC2D2AD3CE2B58C6D68CCC0485DA4FF09A8AE8F5007CB";
   constant CPIX_NORMAL_INIT_37_BIT_01_C : bit_vector(255 downto 0) := x"87DBB10AB2B3DF2DD6A6B80F30D5579BF59BA71B312ACE3C1D5C79227DDD3D50";
   constant CPIX_NORMAL_INIT_37_BIT_02_C : bit_vector(255 downto 0) := x"203ECDB11395E1929E0F26267E5535FE540A359D2C942E6116BC60AE1265BAA0";
   constant CPIX_NORMAL_INIT_37_BIT_03_C : bit_vector(255 downto 0) := x"FBC653543B4EF20C9F48CE8F9D617277657292B9AAAF6CF08E6FEF727428EF6D";
   constant CPIX_NORMAL_INIT_37_BIT_04_C : bit_vector(255 downto 0) := x"7740AF6E886506CF898CB250BD75F268CC4C7253AA0F6A61508A0DE6FA178DB8";
   constant CPIX_NORMAL_INIT_37_BIT_05_C : bit_vector(255 downto 0) := x"292FBB97C5672C495385DB24AC6873CB416B0723C99369849FA94BB4D66E64D2";
   constant CPIX_NORMAL_INIT_37_BIT_06_C : bit_vector(255 downto 0) := x"0276D3276FC010BB7EADB317C149C30ADBC6084A023D63FC5785FD91D96EBDF3";
   constant CPIX_NORMAL_INIT_37_BIT_07_C : bit_vector(255 downto 0) := x"332C319D8553E5A0C8D664351B684AEF8EFD3C01978ADEF3B15A4597B7191229";
   constant CPIX_NORMAL_INIT_37_BIT_08_C : bit_vector(255 downto 0) := x"652435A38FE1432424FA4362FD6E85BC8D19C4A80D5E54DB6A5B9440794C21C6";
   constant CPIX_NORMAL_INIT_37_BIT_09_C : bit_vector(255 downto 0) := x"1347068B930AE7974986C270FB57E019A904B60E62E37A1CCABE2C0B2CE25FDF";
   constant CPIX_NORMAL_INIT_37_BIT_10_C : bit_vector(255 downto 0) := x"9C36BD8292B8EFA2BF1DC1C7C8385DE3C9019129DBACA89660CA782EBE2C3626";
   constant CPIX_NORMAL_INIT_37_BIT_11_C : bit_vector(255 downto 0) := x"0C633C0EEF958334463B937F17B05226A779B114F6A539EBCC844AAB37173EF6";
   constant CPIX_NORMAL_INIT_37_BIT_12_C : bit_vector(255 downto 0) := x"2CE890097B537B7889BDB93FAE2262E558173432E9A35067372B691D0B3CA11C";
   constant CPIX_NORMAL_INIT_37_BIT_13_C : bit_vector(255 downto 0) := x"090D7FD227277C2ADC2D2E58D271A67880738CAB2F9933479FCDCB2BA2EABF5A";
   constant CPIX_NORMAL_INIT_37_BIT_14_C : bit_vector(255 downto 0) := x"3063E590E9545AED959EAF955ACB9E23855072F5515664A498F874FCCF4B48F4";
   constant CPIX_NORMAL_INIT_38_BIT_00_C : bit_vector(255 downto 0) := x"1917D4DED921B1FB746A3F533FF797F4E76F466ECD43A2C0607A34A6E04C7023";
   constant CPIX_NORMAL_INIT_38_BIT_01_C : bit_vector(255 downto 0) := x"D06A4938E5E4D83DFA0F963CBB586CC2FFAD23C3C936A9A512B66CFB58CCEB61";
   constant CPIX_NORMAL_INIT_38_BIT_02_C : bit_vector(255 downto 0) := x"1FE54E80767FC157F4A82C662CB36093842AC8183ACF9944914DECAE2C32B7CC";
   constant CPIX_NORMAL_INIT_38_BIT_03_C : bit_vector(255 downto 0) := x"B39D9601194E04AAE1775C00D5D5816DE667C375C0FDB2E73C3DCDEB7F16AA97";
   constant CPIX_NORMAL_INIT_38_BIT_04_C : bit_vector(255 downto 0) := x"87B68D50E5422DEB12E2586550B71CAE67493FCA21A686F5C6783D14E7428371";
   constant CPIX_NORMAL_INIT_38_BIT_05_C : bit_vector(255 downto 0) := x"05A6D9E3604444809B350FCBB6F5F4F2C325D6EBAD2E399A6F3FD8CD4BFAFC01";
   constant CPIX_NORMAL_INIT_38_BIT_06_C : bit_vector(255 downto 0) := x"966EDB52966111974A4C247906540ED0FE91EDBE9DCDF3AE9F1FBCB5B2302CC5";
   constant CPIX_NORMAL_INIT_38_BIT_07_C : bit_vector(255 downto 0) := x"96734CF040158D07A9F039B5A769701F592B93956372AF13997085D224496B57";
   constant CPIX_NORMAL_INIT_38_BIT_08_C : bit_vector(255 downto 0) := x"F94F340AFE01CAC60A55C22A34EC5B8372588718F98000B447D42BDB31446549";
   constant CPIX_NORMAL_INIT_38_BIT_09_C : bit_vector(255 downto 0) := x"E8F0BD7C5EE42188D7F5A6217A181FA2381FDAE454BE5455BDD5C2A7242D05A7";
   constant CPIX_NORMAL_INIT_38_BIT_10_C : bit_vector(255 downto 0) := x"C738675E7F5DBEF83BF2D600DD5FA2D9B0735F57584EDC907AB1B551034D754A";
   constant CPIX_NORMAL_INIT_38_BIT_11_C : bit_vector(255 downto 0) := x"73BB0C4F8A1E469CCB984BB7BBADB59F6203756F6ECE950986E78C4EFB455CE8";
   constant CPIX_NORMAL_INIT_38_BIT_12_C : bit_vector(255 downto 0) := x"0220D8CAFF9BB7DFE0B18DF756DE48429E4A8C613A11FA7E3B73C94DF6D600D8";
   constant CPIX_NORMAL_INIT_38_BIT_13_C : bit_vector(255 downto 0) := x"D5808E792873F5AACE442EDAA68AA56006796C3C459FB4BF989C42E76C5AF730";
   constant CPIX_NORMAL_INIT_38_BIT_14_C : bit_vector(255 downto 0) := x"677F8089DE151E56FACF6923B7E89C2422E6C982B4C0CBD32F2D14B6FAF6E3E2";
   constant CPIX_NORMAL_INIT_39_BIT_00_C : bit_vector(255 downto 0) := x"79008293BAD3C998A546B6BD484F2FDA338E40DF43172F2F790FF206DBF3404E";
   constant CPIX_NORMAL_INIT_39_BIT_01_C : bit_vector(255 downto 0) := x"0300B9AF4DA65B870E81C4F89C0BE4D39250D599C7A7C47BC1EDAFACB263873C";
   constant CPIX_NORMAL_INIT_39_BIT_02_C : bit_vector(255 downto 0) := x"37DC17E9D5D8F94C84869FC9F84B197EE6D1601C14F3799E58633018607BE12A";
   constant CPIX_NORMAL_INIT_39_BIT_03_C : bit_vector(255 downto 0) := x"4D2941FC4CA3D8C9D396A775701AD4050DC0D90ADE279F25A63D8ADEAC97E289";
   constant CPIX_NORMAL_INIT_39_BIT_04_C : bit_vector(255 downto 0) := x"F957CB9FD035BE823CEA2070580C5DF06AE5D5CB570469ACF7D5FAF00A0E5132";
   constant CPIX_NORMAL_INIT_39_BIT_05_C : bit_vector(255 downto 0) := x"CC82E2FCDDC46695D5692C71B873AB869287F8199E92EC179798788FE0FF47A0";
   constant CPIX_NORMAL_INIT_39_BIT_06_C : bit_vector(255 downto 0) := x"434DBB7F303D84AF2742CB28EEBE4266D765D7CDA61EE11F54711D44A8A0519F";
   constant CPIX_NORMAL_INIT_39_BIT_07_C : bit_vector(255 downto 0) := x"7DDB3E946AB1FBB5E8CCA2668FB3BC0AF0C72BBB1965811627703265EBE7F7AC";
   constant CPIX_NORMAL_INIT_39_BIT_08_C : bit_vector(255 downto 0) := x"9BCC64B824C9F60381BD61D5E7792635F4ABDA7FF067BBA83B6DE213423A1323";
   constant CPIX_NORMAL_INIT_39_BIT_09_C : bit_vector(255 downto 0) := x"349DC358553A1DE05E924795FD56ACF149EB76438CD5A242BBC8D8FAEDAA7605";
   constant CPIX_NORMAL_INIT_39_BIT_10_C : bit_vector(255 downto 0) := x"6AC7152273190AD3C7451AAA4C2247299A97B7B4B4CB4202AB5BBD8B1F3E4E49";
   constant CPIX_NORMAL_INIT_39_BIT_11_C : bit_vector(255 downto 0) := x"F5448A19C47D03188D31987AA82DCA0833FE9A1B265ADD520E70659017C2B6CF";
   constant CPIX_NORMAL_INIT_39_BIT_12_C : bit_vector(255 downto 0) := x"7B220476C9D406447BCA84882C3294A4123786C8B433B3FDAA1BA975D7AF4A97";
   constant CPIX_NORMAL_INIT_39_BIT_13_C : bit_vector(255 downto 0) := x"C56A32AE379EFC7DF5A43A091D57F3BF5E553BC07F82269CE2790C392D529F4E";
   constant CPIX_NORMAL_INIT_39_BIT_14_C : bit_vector(255 downto 0) := x"9F9A68742FFAF821AE05779DE49033991954FEDE1067030A66BE5C2CE754D130";
   constant CPIX_NORMAL_INIT_3A_BIT_00_C : bit_vector(255 downto 0) := x"73FBDD3E55AF85BFDE72B4B5492ECF5DDC107DC180A3661B1BD5895EC74A16E6";
   constant CPIX_NORMAL_INIT_3A_BIT_01_C : bit_vector(255 downto 0) := x"81829A51C45CF5A8179B22864DCEF36419CC0C13DC7EF1A3EAE5D50121A5BDE7";
   constant CPIX_NORMAL_INIT_3A_BIT_02_C : bit_vector(255 downto 0) := x"743CE22EBCBE1AED6CBEAC87970E1E61CC5F15CD5119E8D6D79E909E25A5A8AC";
   constant CPIX_NORMAL_INIT_3A_BIT_03_C : bit_vector(255 downto 0) := x"BCBA48723C51EEC31621A61906276E94981535E0F3909EC2BD3489AD4AC93863";
   constant CPIX_NORMAL_INIT_3A_BIT_04_C : bit_vector(255 downto 0) := x"E748BA597EB895A160D1384254F5FD777BCF442BB98E7539420F6BE1F8A13885";
   constant CPIX_NORMAL_INIT_3A_BIT_05_C : bit_vector(255 downto 0) := x"2F9CA4D39FBA384C17A01A458B38DDD722C40409F2BB33B7176804225ACFDA88";
   constant CPIX_NORMAL_INIT_3A_BIT_06_C : bit_vector(255 downto 0) := x"32115B52C96BD7C23238A49574E673271B0D2C482F0274CE2FCD0C847DB4AAB2";
   constant CPIX_NORMAL_INIT_3A_BIT_07_C : bit_vector(255 downto 0) := x"BE923026FACE8D140FA1A3F21E4225783C84C8CD86578C6A160CD57FC0636DC7";
   constant CPIX_NORMAL_INIT_3A_BIT_08_C : bit_vector(255 downto 0) := x"081AB243F667F947A23ED28CBEA787C931E4E2AE416ED2E00FA58875D488BF97";
   constant CPIX_NORMAL_INIT_3A_BIT_09_C : bit_vector(255 downto 0) := x"8947DFD0CBBAD6A206556F932B3B2D273A0CFC9705F00F4320C039063F16DA49";
   constant CPIX_NORMAL_INIT_3A_BIT_10_C : bit_vector(255 downto 0) := x"1E461B9D25D1DEED858ACCA00C776963ADE265095F93C95984B9038F3B942DF2";
   constant CPIX_NORMAL_INIT_3A_BIT_11_C : bit_vector(255 downto 0) := x"6C059D15DBA726595F503C4A4B246B348151AF9DB6E1F16D27768DC9576B669E";
   constant CPIX_NORMAL_INIT_3A_BIT_12_C : bit_vector(255 downto 0) := x"8E3FAD98BDA1E29ED559073AF1FA36BC508D4907F0D831F2CA3445EAF1545F5E";
   constant CPIX_NORMAL_INIT_3A_BIT_13_C : bit_vector(255 downto 0) := x"20432FF2AFCFDF05D4C0407E5F41E886324034350B78658FF1BDF379D35457A7";
   constant CPIX_NORMAL_INIT_3A_BIT_14_C : bit_vector(255 downto 0) := x"9AA43B94B3EA303D70E67996D0267583AA36A72AB3D7D0C9EE73F74041D58970";
   constant CPIX_NORMAL_INIT_3B_BIT_00_C : bit_vector(255 downto 0) := x"43CDCDFDF9492F8FE78A894F2B435FFADCE3430F4034E68F117A14A77B58B4BC";
   constant CPIX_NORMAL_INIT_3B_BIT_01_C : bit_vector(255 downto 0) := x"8D32EBB0C8CDF689210063A9059AA347820B54AEE9BBA9AAB820FF98EE0268A3";
   constant CPIX_NORMAL_INIT_3B_BIT_02_C : bit_vector(255 downto 0) := x"5E8384195DC00B75CC35EE2F08554BC6FCED4B655CA95EBA387FE3324A514439";
   constant CPIX_NORMAL_INIT_3B_BIT_03_C : bit_vector(255 downto 0) := x"ABDA3FFC9B12930D02CF9E7C5CD160321770175771D40C7E5A4BD733596CBA18";
   constant CPIX_NORMAL_INIT_3B_BIT_04_C : bit_vector(255 downto 0) := x"5F1378419D809270512741A8859D3CD9E3B4A42C03CAB5A9E606C010057A469A";
   constant CPIX_NORMAL_INIT_3B_BIT_05_C : bit_vector(255 downto 0) := x"0351B1A10955C96FB12655A26E13674633A3B00241C4F485B3B394042AC8FCC0";
   constant CPIX_NORMAL_INIT_3B_BIT_06_C : bit_vector(255 downto 0) := x"552A5974EC89F50C4EF57278C9DDEF21A2F3D0583678DA62131C40194F098D7F";
   constant CPIX_NORMAL_INIT_3B_BIT_07_C : bit_vector(255 downto 0) := x"0F550A58445D3F40FC5727578CBFCA2F2BB8BCC7F53CD1F09019702831E2C14E";
   constant CPIX_NORMAL_INIT_3B_BIT_08_C : bit_vector(255 downto 0) := x"BD43D862B70C5ABECA7A71B4A6799A8F2E1F1AF8694E21581EE2DD627DF882B2";
   constant CPIX_NORMAL_INIT_3B_BIT_09_C : bit_vector(255 downto 0) := x"8F714E506DE960FFFB58C83953EDE8588623CFE458A77FD3097152A98DB53D22";
   constant CPIX_NORMAL_INIT_3B_BIT_10_C : bit_vector(255 downto 0) := x"B744D002A4132144913BB39198287BE705089A844A6A4A6582CA3C20B7C33B47";
   constant CPIX_NORMAL_INIT_3B_BIT_11_C : bit_vector(255 downto 0) := x"8423BF3351BD667F195D1CBEA4BB406F84915ED78220B3440173087683258160";
   constant CPIX_NORMAL_INIT_3B_BIT_12_C : bit_vector(255 downto 0) := x"0B15A09CAF996ABA0B630A37785457DFB110AF7E91CFD02AB9A0D7870AD9ADF1";
   constant CPIX_NORMAL_INIT_3B_BIT_13_C : bit_vector(255 downto 0) := x"1DCB9A80B8A288EA9A44EEA692CB6D86479BD872B5AD612B7D93FFD3E49827AC";
   constant CPIX_NORMAL_INIT_3B_BIT_14_C : bit_vector(255 downto 0) := x"0F934032C83D51FE12AC283F60E29AB3B2EFB43CC3F22CA04CF4E7DF510F63AF";
   constant CPIX_NORMAL_INIT_3C_BIT_00_C : bit_vector(255 downto 0) := x"18A4D0854342B430C46EF262FAC30EF46ACB32BF0DA4F22D1A4E485B0FC3444B";
   constant CPIX_NORMAL_INIT_3C_BIT_01_C : bit_vector(255 downto 0) := x"C2FCCEE3017A06F1E2BA70FD9B5FE799916EB831263BFE9185C5DBBC690348FD";
   constant CPIX_NORMAL_INIT_3C_BIT_02_C : bit_vector(255 downto 0) := x"EF563843906B1456B6125468A6A139BBDDF4D23A4238E7B0FA4D99A021D8B12E";
   constant CPIX_NORMAL_INIT_3C_BIT_03_C : bit_vector(255 downto 0) := x"57C1D4B220880B6673705DB4E38F612322AE1BC22857A6F40DEFE2AAA6137995";
   constant CPIX_NORMAL_INIT_3C_BIT_04_C : bit_vector(255 downto 0) := x"1F48DFA97810EB577B1AA69C82857B4914A69A6B49E37DF053BFA8C6DE1C2DD1";
   constant CPIX_NORMAL_INIT_3C_BIT_05_C : bit_vector(255 downto 0) := x"64E186FE42BBB3195352372A45E37BCD71A553EB186875973FE544EAF4E94C75";
   constant CPIX_NORMAL_INIT_3C_BIT_06_C : bit_vector(255 downto 0) := x"46C623518D76E8472A1A7142741B2B7F573786B5B899F7868873F0731513B60B";
   constant CPIX_NORMAL_INIT_3C_BIT_07_C : bit_vector(255 downto 0) := x"5302389714C8C76D0AE9DDE10ED8B243638FA17A6D91B5B3DE8D9C3B8E8E16AD";
   constant CPIX_NORMAL_INIT_3C_BIT_08_C : bit_vector(255 downto 0) := x"16A7FCEF5DBD09543BE17F1BACC7EF835ED262B0FB45814E96431DFF6C5690AA";
   constant CPIX_NORMAL_INIT_3C_BIT_09_C : bit_vector(255 downto 0) := x"3C8F85557668F7AC4302900E23ACFD1704CDF742334A80E0F270D2F4F5F092ED";
   constant CPIX_NORMAL_INIT_3C_BIT_10_C : bit_vector(255 downto 0) := x"1C3699A81EE0911901347706B7B1C0C8200798D465A650952627FD534280848F";
   constant CPIX_NORMAL_INIT_3C_BIT_11_C : bit_vector(255 downto 0) := x"D82B4267B844548E6EB9CFFE41F37BA103AE684528C11EE03A5A8C79ABFC7669";
   constant CPIX_NORMAL_INIT_3C_BIT_12_C : bit_vector(255 downto 0) := x"1E19CF6BE75E26BB9AD8BE83C3C2BC3262DD84B313E9AD433464AF8273544B24";
   constant CPIX_NORMAL_INIT_3C_BIT_13_C : bit_vector(255 downto 0) := x"44CCB8BDB0018E8BEBF7AD8732384A86A7C3E47BC35CF72A184DFDB755D111BA";
   constant CPIX_NORMAL_INIT_3C_BIT_14_C : bit_vector(255 downto 0) := x"19064AD78C2AFFC2D68F32A06FB364454D5B51C5AC74EFC8097017C09AD2862C";
   constant CPIX_NORMAL_INIT_3D_BIT_00_C : bit_vector(255 downto 0) := x"0FDA4C586363B47603F87318518370E91323BE56379DB22F3B51D4114F0C70DD";
   constant CPIX_NORMAL_INIT_3D_BIT_01_C : bit_vector(255 downto 0) := x"D0560EEF8835C8A5555AA60003852C91157838E851879A9618F1FE7959803DF1";
   constant CPIX_NORMAL_INIT_3D_BIT_02_C : bit_vector(255 downto 0) := x"4BDF499BC05A32013C17EC17AB6A49ABEC9579B7DEFF98F305C6C6EE6ED213EC";
   constant CPIX_NORMAL_INIT_3D_BIT_03_C : bit_vector(255 downto 0) := x"90F02168D2AB6B0FCA95C1C9987F368CCCE54DF1FE25F07A2E0229ABBC798035";
   constant CPIX_NORMAL_INIT_3D_BIT_04_C : bit_vector(255 downto 0) := x"21CA3A9C6335BD25143859CB53AFDA1B1F61F4BF1B1A80223A15E29D1B07CDB0";
   constant CPIX_NORMAL_INIT_3D_BIT_05_C : bit_vector(255 downto 0) := x"941FE1173530EFDE370AF83A4486883CB79E83E6AC31195E00A92572D30F78F8";
   constant CPIX_NORMAL_INIT_3D_BIT_06_C : bit_vector(255 downto 0) := x"A8FD2D66FEF41D889682F74B0EB7A1F7C4596D1D4AB85B3D98F9339C1325FE6F";
   constant CPIX_NORMAL_INIT_3D_BIT_07_C : bit_vector(255 downto 0) := x"F706DB60172B419176E6B9EF388777B3B02776C048B427C37363EEED992CDBCF";
   constant CPIX_NORMAL_INIT_3D_BIT_08_C : bit_vector(255 downto 0) := x"3958C4B8E24CEA716C25345ECCD19E6BC21D0B0360A8778C1A5495DAC1810CB3";
   constant CPIX_NORMAL_INIT_3D_BIT_09_C : bit_vector(255 downto 0) := x"4B95315AFEE9AB0E75D3D8531B05C4F05EC78A5A48688DABAB6D3516981072C1";
   constant CPIX_NORMAL_INIT_3D_BIT_10_C : bit_vector(255 downto 0) := x"DD4A1736947C15AD723B805C45046B2746AE9392289A6266770F43BBFADFEE5D";
   constant CPIX_NORMAL_INIT_3D_BIT_11_C : bit_vector(255 downto 0) := x"E83522F95815166912084D8E468B16D6C4FA209CF8DA1CEDB3646F771E1C1C76";
   constant CPIX_NORMAL_INIT_3D_BIT_12_C : bit_vector(255 downto 0) := x"F4C80881564B019656E19F7F46F7016614E9DE26CF90B8E6C3E9949EF7BF9544";
   constant CPIX_NORMAL_INIT_3D_BIT_13_C : bit_vector(255 downto 0) := x"A456DA1E3E77504BC2783C88F51C71AE02584F38D64F8D13989C601D565B120B";
   constant CPIX_NORMAL_INIT_3D_BIT_14_C : bit_vector(255 downto 0) := x"37C0D0DCC336EB2DCF5AA28D0C14DF824D01B78BDFC50F7CDD6018DF9A8E01FC";
   constant CPIX_NORMAL_INIT_3E_BIT_00_C : bit_vector(255 downto 0) := x"E6DCBD7B2A333B26E34F7B53C688B04BDB70B3C1474D7D59DCE93EDD1B346D63";
   constant CPIX_NORMAL_INIT_3E_BIT_01_C : bit_vector(255 downto 0) := x"92CE4154EBF10F8C35E71F8C7F581D67065D531C09585044851B9206FEAA8F1F";
   constant CPIX_NORMAL_INIT_3E_BIT_02_C : bit_vector(255 downto 0) := x"F7830C73557E405ED053ECB0826AC45BFBE01BDD67740F2A7C2DF4F58667A734";
   constant CPIX_NORMAL_INIT_3E_BIT_03_C : bit_vector(255 downto 0) := x"A96B3E90ED603BC73555FB2D5EC837D499EAC24DC2E3F58C99B148F385347043";
   constant CPIX_NORMAL_INIT_3E_BIT_04_C : bit_vector(255 downto 0) := x"CF8001FDF64934E9587E8CE04A30EBB5CF84FFCBD3B634D9FF4D68891594A4EF";
   constant CPIX_NORMAL_INIT_3E_BIT_05_C : bit_vector(255 downto 0) := x"0E5D638953FF506F29A6161B5A1A4ED7A041C5A06F6452A9991E728177094A54";
   constant CPIX_NORMAL_INIT_3E_BIT_06_C : bit_vector(255 downto 0) := x"83A4DD4094BDF47D16C5402A191F41FB02387BD46BDB7B7A9CB30FEDCE1A7CB5";
   constant CPIX_NORMAL_INIT_3E_BIT_07_C : bit_vector(255 downto 0) := x"A622A99A03AEA19D997F091DFB7B26A54C8E24C07BB7C9EE55F3E7A32020B00B";
   constant CPIX_NORMAL_INIT_3E_BIT_08_C : bit_vector(255 downto 0) := x"0FFB3B7A5D25F6EF04FE0588F081C30F8A24E9D0E268278EC89A1428C8E58392";
   constant CPIX_NORMAL_INIT_3E_BIT_09_C : bit_vector(255 downto 0) := x"5FA9E8DE692B0C0DC2C309CB64C1E4B99D95355050A66EFDE7A38326D1156624";
   constant CPIX_NORMAL_INIT_3E_BIT_10_C : bit_vector(255 downto 0) := x"1C5322CE6391EC494CAB0D04ED221B218D07CC109FBDA736C691FC080A7A2E9B";
   constant CPIX_NORMAL_INIT_3E_BIT_11_C : bit_vector(255 downto 0) := x"94E48D83A766BF7556F9C0D551CED855871019931ACAFEC700180F3C9AFE4361";
   constant CPIX_NORMAL_INIT_3E_BIT_12_C : bit_vector(255 downto 0) := x"12FD479DA54B5596480DB88621A907B5014F5D0DEF8B0FF581FF2CEC8400119B";
   constant CPIX_NORMAL_INIT_3E_BIT_13_C : bit_vector(255 downto 0) := x"8973152342047DE5186B27AAAA5FC6AC025C36BF8636CA13821AED1B5EB29E89";
   constant CPIX_NORMAL_INIT_3E_BIT_14_C : bit_vector(255 downto 0) := x"3CA4F559F7A8413F328E08875A9DA9B8B03F3AAF1DD01FCBB635B508AE758B8E";
   constant CPIX_NORMAL_INIT_3F_BIT_00_C : bit_vector(255 downto 0) := x"4F0176ED501A42A4DD38CB8E51F6CB674D580D43C517A4041359BBE2A9B98962";
   constant CPIX_NORMAL_INIT_3F_BIT_01_C : bit_vector(255 downto 0) := x"93F05E06021CFCBB01E5A0E85587ECFBB8B17A2CEFD557C281B87883A55ADC0A";
   constant CPIX_NORMAL_INIT_3F_BIT_02_C : bit_vector(255 downto 0) := x"FE77EDB9E447A72FFEB7531AB2AD5A47F3B0B45C1C65C343EA4F82C9FC9434BA";
   constant CPIX_NORMAL_INIT_3F_BIT_03_C : bit_vector(255 downto 0) := x"FFF7DEEFB6737C5FDE1CAF465DBFF86A35B3E9652AAA9F5B6E776F8AF2A651F4";
   constant CPIX_NORMAL_INIT_3F_BIT_04_C : bit_vector(255 downto 0) := x"530EA4FD10962CDD118778D07333AD734644BC38D4062E60613604AF3F05D6F3";
   constant CPIX_NORMAL_INIT_3F_BIT_05_C : bit_vector(255 downto 0) := x"3329FE835FA92A1D01F01433369ED64F06093DF43482EF531C089BBD90F7354E";
   constant CPIX_NORMAL_INIT_3F_BIT_06_C : bit_vector(255 downto 0) := x"12A1C0D358BAB56B33BD5CC6326C1D4B0486CA848268172B0950A79B1BFEA407";
   constant CPIX_NORMAL_INIT_3F_BIT_07_C : bit_vector(255 downto 0) := x"12284D875B80F48F5350FC6AB4D568509988B5664033E3EA3E30497E3D35734F";
   constant CPIX_NORMAL_INIT_3F_BIT_08_C : bit_vector(255 downto 0) := x"0A6C2F2108C793FF3379DFF10824FB6218816DD5990502110F18AC2BA8FB76FE";
   constant CPIX_NORMAL_INIT_3F_BIT_09_C : bit_vector(255 downto 0) := x"024189369B8B56AD2245AA5B58FCB4563B8ADB42AA4C2E6D85B0C3A0F438DF7C";
   constant CPIX_NORMAL_INIT_3F_BIT_10_C : bit_vector(255 downto 0) := x"0453D0BE1EDF6A4920B2B5750A77DE7A3C096E7F163CD22D95083049E3B94DAA";
   constant CPIX_NORMAL_INIT_3F_BIT_11_C : bit_vector(255 downto 0) := x"0251E03A740FE329210765F83902BF042222DD961FE4381083A19A926CEF35CB";
   constant CPIX_NORMAL_INIT_3F_BIT_12_C : bit_vector(255 downto 0) := x"0219C5080596F28314C47F1806E27A582C3A3B3D003259F198032B70640AABF6";
   constant CPIX_NORMAL_INIT_3F_BIT_13_C : bit_vector(255 downto 0) := x"0210690A5C80A3E50A6141D12E2F08D40A7E964D973FF615145C89B588EA24E1";
   constant CPIX_NORMAL_INIT_3F_BIT_14_C : bit_vector(255 downto 0) := x"0008251613988182B046C4C19AF065CC4E76358A5A15606F4D207336E170E24A";
   constant CPIX_NORMAL_INIT_40_BIT_00_C : bit_vector(255 downto 0) := x"3404839B7E4C094A6E410BB957459E384D57B7D68C3E8A494DEA433D79BB36D2";
   constant CPIX_NORMAL_INIT_40_BIT_01_C : bit_vector(255 downto 0) := x"C67B45817359CF5FB7B9CA199A38CB7BE1FEED8415DAA0E79BC46BE88C3F55EB";
   constant CPIX_NORMAL_INIT_40_BIT_02_C : bit_vector(255 downto 0) := x"EC68B6BE841BE303D8ED5EABCADE1B43F19BA4C3B95B54A5FF070875CE3D7BEB";
   constant CPIX_NORMAL_INIT_40_BIT_03_C : bit_vector(255 downto 0) := x"758E7589912EE80A33E2E40DA51BA85765E1367C8FC2F4FC9A9D407846FA1DEB";
   constant CPIX_NORMAL_INIT_40_BIT_04_C : bit_vector(255 downto 0) := x"4E0FB6006D1AFE8D07CFB2B550450A7275A4AFF4C710F3BFD27D1D9BF04734ED";
   constant CPIX_NORMAL_INIT_40_BIT_05_C : bit_vector(255 downto 0) := x"543B3AF6FBB6E84D39E9288BA833ABD3756E59FE888AC9A5F11785874173E19F";
   constant CPIX_NORMAL_INIT_40_BIT_06_C : bit_vector(255 downto 0) := x"6D80F87B57E26CA31635FB9CF7D7F10678212D21BF29A725BB9F3557D7B8A7EF";
   constant CPIX_NORMAL_INIT_40_BIT_07_C : bit_vector(255 downto 0) := x"00115B54B76E52F2A76C64C0FFD0411A41EBEC40FAB63E6B32CED3AAF13B9DDF";
   constant CPIX_NORMAL_INIT_40_BIT_08_C : bit_vector(255 downto 0) := x"37D6DD6AC03761D8975A0761C01CF34751880A23D7DE543D72EBF5405DF7705D";
   constant CPIX_NORMAL_INIT_40_BIT_09_C : bit_vector(255 downto 0) := x"B1910870C17B75A5E545C8238DFC62293587509542DFA16858B54FD2757E3EAD";
   constant CPIX_NORMAL_INIT_40_BIT_10_C : bit_vector(255 downto 0) := x"1694D024F4647878831B57D43B4D922950FC885EE358403B57EB97E45FB48FA1";
   constant CPIX_NORMAL_INIT_40_BIT_11_C : bit_vector(255 downto 0) := x"09297ACDADA3CBFE025CA0D715AF370D440B52CEDDBA17457CD879028C75C6A5";
   constant CPIX_NORMAL_INIT_40_BIT_12_C : bit_vector(255 downto 0) := x"0B3CAFB9616C1D302FD82709F5ECB8B05676B340C4C57223191ED3CC2F27A035";
   constant CPIX_NORMAL_INIT_40_BIT_13_C : bit_vector(255 downto 0) := x"366AF9045E5D65F20639114E0E254F941EBFCA7F15E83B9A00A01A7C91E5F405";
   constant CPIX_NORMAL_INIT_40_BIT_14_C : bit_vector(255 downto 0) := x"59BBAE5F9B511D164A1B3DED33BE5D739E1ACC26E295EE484CA9E9C723016E11";
   constant CPIX_NORMAL_INIT_41_BIT_00_C : bit_vector(255 downto 0) := x"C867B11B5A0D1D2B8DD434E39488A1992A8937B7CA4769697338E4585BB476BD";
   constant CPIX_NORMAL_INIT_41_BIT_01_C : bit_vector(255 downto 0) := x"B964D7858CDAA24E61D4B81EC6700FBCF9151B34C1482D3F4B35F81082A71C97";
   constant CPIX_NORMAL_INIT_41_BIT_02_C : bit_vector(255 downto 0) := x"B9A848F155509EBA3FF66A8CB6E4AF6BBF35231C57E3A337C21874CA20C2D5CD";
   constant CPIX_NORMAL_INIT_41_BIT_03_C : bit_vector(255 downto 0) := x"05C0FC773E3EE12554790BFBD1D0E3E94DC48BE06632D578E688E71045CC87AE";
   constant CPIX_NORMAL_INIT_41_BIT_04_C : bit_vector(255 downto 0) := x"98F9879B52C84AA5A5CA4CD9C1BD2011F20A4C1F6557A20909A00FFF2D5A4E61";
   constant CPIX_NORMAL_INIT_41_BIT_05_C : bit_vector(255 downto 0) := x"96C878D1DF999CBBA4029FEE932E0D0E1BFEE3CDA4BF27E7AFFEF632AA6D4189";
   constant CPIX_NORMAL_INIT_41_BIT_06_C : bit_vector(255 downto 0) := x"CB00315E4D69ECAEB714D0AE125AFAB9BC65ED3E0228E4E05F22782816E9228D";
   constant CPIX_NORMAL_INIT_41_BIT_07_C : bit_vector(255 downto 0) := x"6CC7A36E1D66756E40FDBDDB9BA4C163FDD167241D7E363F18CB449C01B55F07";
   constant CPIX_NORMAL_INIT_41_BIT_08_C : bit_vector(255 downto 0) := x"7259D29593FF4E481A9B17A9C11E343587442CA3DE531FAF793EF5A9BB80DD6F";
   constant CPIX_NORMAL_INIT_41_BIT_09_C : bit_vector(255 downto 0) := x"BB927CFF38C996AA780AC18B907916AE098F0196E3F78BC7AC13FE54C05F2A3B";
   constant CPIX_NORMAL_INIT_41_BIT_10_C : bit_vector(255 downto 0) := x"B44E29DBA8640A76EC74DA3F57C4275C4C838B488139F66C220E816F1133314B";
   constant CPIX_NORMAL_INIT_41_BIT_11_C : bit_vector(255 downto 0) := x"DAF40022858EBD1668EC1E16D7FA4BD92DA011A07BFE1296D3DDF1E0581A8C72";
   constant CPIX_NORMAL_INIT_41_BIT_12_C : bit_vector(255 downto 0) := x"C1202FBE8FC03EEEA11B287FB3C39CFACB6974F6EA4475CA132F5685EE7CB43E";
   constant CPIX_NORMAL_INIT_41_BIT_13_C : bit_vector(255 downto 0) := x"4E1784EEEA5251D51B3004BE8C29B29465F9E495A352FFB2FF299D56403D5B98";
   constant CPIX_NORMAL_INIT_41_BIT_14_C : bit_vector(255 downto 0) := x"6193F8451A0F499DB0B22B17B9DC6528B6A2F1C9175D21C08D46C86C148F9F02";
   constant CPIX_NORMAL_INIT_42_BIT_00_C : bit_vector(255 downto 0) := x"C164989C8030892539B53B6E4B7A7302924F83DB486F33CD9380884FA8EEF8FD";
   constant CPIX_NORMAL_INIT_42_BIT_01_C : bit_vector(255 downto 0) := x"BACBFDAA0D477CEDC9B234030AE4E9826F8BFA49F3CDB5C37DA6B08BEA377A06";
   constant CPIX_NORMAL_INIT_42_BIT_02_C : bit_vector(255 downto 0) := x"3D1CACBF25A85E492E11A9D8E9829624C320FBCEC2410AD20DE67983B693249E";
   constant CPIX_NORMAL_INIT_42_BIT_03_C : bit_vector(255 downto 0) := x"6B2F07D2F9F190F35AB11F0E9FE6AAB431033C4F5B255F5DAFF48E2294B3AA78";
   constant CPIX_NORMAL_INIT_42_BIT_04_C : bit_vector(255 downto 0) := x"D0768A7672A567397DBD9D7292138A0A265406D1E7AD2C70AA364CFD74F0415C";
   constant CPIX_NORMAL_INIT_42_BIT_05_C : bit_vector(255 downto 0) := x"FD950BF63B6E525E83064DA6EE000F672B77D8DE2CE1F14F0ADE310ECDDC8B55";
   constant CPIX_NORMAL_INIT_42_BIT_06_C : bit_vector(255 downto 0) := x"DC9325993AA8008C3F6F5465BB57F52D8AFBEECD719318AA6E438C510EA97EE0";
   constant CPIX_NORMAL_INIT_42_BIT_07_C : bit_vector(255 downto 0) := x"D6D83C3050127BC9338DFA98642D2B72CF342E22DDDE48CCD3C7546DD7E75BFA";
   constant CPIX_NORMAL_INIT_42_BIT_08_C : bit_vector(255 downto 0) := x"2C0A9D3F592684ACAAB0E082F1402296C7F771E386E6C6F629A24AFD45AFC3D7";
   constant CPIX_NORMAL_INIT_42_BIT_09_C : bit_vector(255 downto 0) := x"D3DB61DEC24E40E77B652D788FAA9932B7AE44A9F5AE9797972E538BA24AA27A";
   constant CPIX_NORMAL_INIT_42_BIT_10_C : bit_vector(255 downto 0) := x"A29C53AEBEB580C6D3ABE4B49C0BBEE31D4F84BB3E3C75B5A854A048E2A424E4";
   constant CPIX_NORMAL_INIT_42_BIT_11_C : bit_vector(255 downto 0) := x"E7B88B15793BBF150D9991A7DD3BEC246F37B69C25BFE3CC32D390718A1412CB";
   constant CPIX_NORMAL_INIT_42_BIT_12_C : bit_vector(255 downto 0) := x"00936F3F8F803F6176B1038F52D7109F0E9D6B6BAD247A35F5190948BB8C0E06";
   constant CPIX_NORMAL_INIT_42_BIT_13_C : bit_vector(255 downto 0) := x"A1FDE5E045C9578D1BE4E298AF7BDAFC9A864B0E769F12F5E936EFAA6FFB4DD9";
   constant CPIX_NORMAL_INIT_42_BIT_14_C : bit_vector(255 downto 0) := x"EE311E2F614BF4B7784AE5C741A5B5C43A9F24E2EA43985C583E63097763DA1F";
   constant CPIX_NORMAL_INIT_43_BIT_00_C : bit_vector(255 downto 0) := x"5606824C8B21C3E2D995B46975C253146D55399E5B31C159699445AF52864109";
   constant CPIX_NORMAL_INIT_43_BIT_01_C : bit_vector(255 downto 0) := x"9FBCBC02537BDD1D76759E9B7D6C21DEAB8223BACD259E43B16F52C82722ACF7";
   constant CPIX_NORMAL_INIT_43_BIT_02_C : bit_vector(255 downto 0) := x"B5787B3B3E00FC695E4FC3A0134F34DA8E921B73499B2FBBD929B80FD7AFDE5A";
   constant CPIX_NORMAL_INIT_43_BIT_03_C : bit_vector(255 downto 0) := x"77DF288793C41AB4946F52D66BC8A6EF0AE2D107B1A2394F063DDB7C5AFD965B";
   constant CPIX_NORMAL_INIT_43_BIT_04_C : bit_vector(255 downto 0) := x"495DFDF4D4455E9D33FE78275A94BFBA128F19EC2E9D0ECB3C7D01152C94AD62";
   constant CPIX_NORMAL_INIT_43_BIT_05_C : bit_vector(255 downto 0) := x"6B3E415402C9FBDE54F5A9B3F3AFF3DC4BBF769BB38A0A151DDBBE401B06EA7E";
   constant CPIX_NORMAL_INIT_43_BIT_06_C : bit_vector(255 downto 0) := x"EDDEA96DBB2C98703AC4161F1043317D3A1FDD84D9CD13BD5E70ECCABC8B1E44";
   constant CPIX_NORMAL_INIT_43_BIT_07_C : bit_vector(255 downto 0) := x"738871FC1F7576BB1296ACC1FAC36C4C5BB6042D8420AC1F2D95628ED509444F";
   constant CPIX_NORMAL_INIT_43_BIT_08_C : bit_vector(255 downto 0) := x"35CB9E5B4237FBC5054F07DBEC9033346B5381D0812F1A6D4207216FCCA34450";
   constant CPIX_NORMAL_INIT_43_BIT_09_C : bit_vector(255 downto 0) := x"3384CFB8A9918297327274689DAE996D5A2934C87EB77C810A2C7C74B74FB3E1";
   constant CPIX_NORMAL_INIT_43_BIT_10_C : bit_vector(255 downto 0) := x"6903682910E66373054A7CAF94E419187738B22E7BC82D782549F4E863FF3BCE";
   constant CPIX_NORMAL_INIT_43_BIT_11_C : bit_vector(255 downto 0) := x"056FCE7247F01FB226C0206500879F29203DE8EFA41C31CCB29AFA44BDBC3A68";
   constant CPIX_NORMAL_INIT_43_BIT_12_C : bit_vector(255 downto 0) := x"3B11D73DDABE1EE4712F73B42D537E0389206793EA9EA545A25C4BD37115733D";
   constant CPIX_NORMAL_INIT_43_BIT_13_C : bit_vector(255 downto 0) := x"340715430508DD87F7AF69196970963C406AEDD4AA6EE27381D0DDAE7D2F77A0";
   constant CPIX_NORMAL_INIT_43_BIT_14_C : bit_vector(255 downto 0) := x"3740AF71C5675E569BBDED32A7484AF75E5D81A7ABC1E0EDCD02E54365727B47";
   constant CPIX_NORMAL_INIT_44_BIT_00_C : bit_vector(255 downto 0) := x"0FBD51B493E000A23210F20478D4671704382C472DD22275569086F78C343AD9";
   constant CPIX_NORMAL_INIT_44_BIT_01_C : bit_vector(255 downto 0) := x"52B9EFCB7FD2FDCA568B21C9B7F7B135A1E1B141117976F42B1DB270BA20B1BD";
   constant CPIX_NORMAL_INIT_44_BIT_02_C : bit_vector(255 downto 0) := x"EA30043E536679F8F39F56551F4863530B75A3BC6D4DC84D64BEEB8794D8749A";
   constant CPIX_NORMAL_INIT_44_BIT_03_C : bit_vector(255 downto 0) := x"4C1C68DEDF22062CD6787F07073F1FA62E386BE672238008CB2999DE5B0A7D6D";
   constant CPIX_NORMAL_INIT_44_BIT_04_C : bit_vector(255 downto 0) := x"16ED40EF673DD1D57683DC21559AEFD51521D2FDDB7A5175A8714D51BC2F7F43";
   constant CPIX_NORMAL_INIT_44_BIT_05_C : bit_vector(255 downto 0) := x"CF101FEB564C0E85D42E1A61557F20B1583D4F0DB08F6607792D78FBD4D22DC2";
   constant CPIX_NORMAL_INIT_44_BIT_06_C : bit_vector(255 downto 0) := x"73F032A7E22FE9C72D69865531E845AB8653A141AC7A9EF4DB0D06CD72924605";
   constant CPIX_NORMAL_INIT_44_BIT_07_C : bit_vector(255 downto 0) := x"8E850E54313C5AEA171CFA1B5D0112FB23585F5A06F351F16701913FEDA87AD9";
   constant CPIX_NORMAL_INIT_44_BIT_08_C : bit_vector(255 downto 0) := x"0282CC5886BB5077DF79FF80883F51C4F0ACC6F9AD35595CDCD502F5B0A1DD2F";
   constant CPIX_NORMAL_INIT_44_BIT_09_C : bit_vector(255 downto 0) := x"A0CE4D0CEC710B746054865D6B360773048446F96CFCBD780D47FC0362366A36";
   constant CPIX_NORMAL_INIT_44_BIT_10_C : bit_vector(255 downto 0) := x"FB1D3399BC2A63DCF37E067C3D4D0F1C6CF4FE6576771EF33A3F118DFB5536EC";
   constant CPIX_NORMAL_INIT_44_BIT_11_C : bit_vector(255 downto 0) := x"2B513F3FF9615EAAEEB1E893BA9CE50E3B82BFCAC5FFA079EC55001D8B2D5C5A";
   constant CPIX_NORMAL_INIT_44_BIT_12_C : bit_vector(255 downto 0) := x"42FF901FD7ECFE269889B1AB7C3C29C5362CF3C69C35A157121C124437F22AE4";
   constant CPIX_NORMAL_INIT_44_BIT_13_C : bit_vector(255 downto 0) := x"6FB64FA4F28819A17D3052A769D4B8B07D15DD41B4AA025942F8EB1370A4B466";
   constant CPIX_NORMAL_INIT_44_BIT_14_C : bit_vector(255 downto 0) := x"EDB52A9D52FF1F1D0ABA2BD55EA501942A87E4EA7B0B2456F3B72D72427C6514";
   constant CPIX_NORMAL_INIT_45_BIT_00_C : bit_vector(255 downto 0) := x"7D018013EC56DD0C3BC657EF072853FE8BEB2362C5817356BB0258A5CF7AE415";
   constant CPIX_NORMAL_INIT_45_BIT_01_C : bit_vector(255 downto 0) := x"B23F8F3DA681156CC814C2BE7BA07E71C12AF15F93EDBFF40DF0231E778105D5";
   constant CPIX_NORMAL_INIT_45_BIT_02_C : bit_vector(255 downto 0) := x"F6F432155FA51CF6EEBF32A2246DAB99CDD192BBB6765969300173ACE9E08688";
   constant CPIX_NORMAL_INIT_45_BIT_03_C : bit_vector(255 downto 0) := x"2300A6BC14A8415A36ECE46FACD9FF7DB61C9CCED6E4C233E5D8EEC7A2EC6983";
   constant CPIX_NORMAL_INIT_45_BIT_04_C : bit_vector(255 downto 0) := x"0B4C5A88C0555A601EECB411105129E713AC90EE23EF63E5925A3E2276CE03FB";
   constant CPIX_NORMAL_INIT_45_BIT_05_C : bit_vector(255 downto 0) := x"B966277CAF750ADFB6B2C60B8408C31807436194C59C183BB9FC86558D747848";
   constant CPIX_NORMAL_INIT_45_BIT_06_C : bit_vector(255 downto 0) := x"74CD6527ECD48B86E5C90F418A3E0535B795D851DC7FD3D481CF8A2E8844A68F";
   constant CPIX_NORMAL_INIT_45_BIT_07_C : bit_vector(255 downto 0) := x"6901B9B74E82D33889A8ADC84640519535E0087DDF63D1E81A318C08C06D93FD";
   constant CPIX_NORMAL_INIT_45_BIT_08_C : bit_vector(255 downto 0) := x"71C236A3FAE54D9086C8014D83BD81DF8B1E55A4A653885726314AE68E022DD3";
   constant CPIX_NORMAL_INIT_45_BIT_09_C : bit_vector(255 downto 0) := x"5908A37B07CB4B9C0D693F5C608D509CBC631EE286582C55B6E5EF67D394D62D";
   constant CPIX_NORMAL_INIT_45_BIT_10_C : bit_vector(255 downto 0) := x"B612C8EEBBC0AA6F9B0FCDED33738FA73D9DA25AE5CE8D54A13615D6F5F53077";
   constant CPIX_NORMAL_INIT_45_BIT_11_C : bit_vector(255 downto 0) := x"1F5C5555ACA42D1DBDB1005B8D206050E2C996E5AA41BA68CB54885B715B9EEE";
   constant CPIX_NORMAL_INIT_45_BIT_12_C : bit_vector(255 downto 0) := x"7C692F30161514C4EC548F794281008D7CA7C5B45CDA954C3CA9095C73195BCD";
   constant CPIX_NORMAL_INIT_45_BIT_13_C : bit_vector(255 downto 0) := x"0CC9F1878A4BF945C51DF54195A81090A354E8B1E85CE8B358C8738A5F54DD23";
   constant CPIX_NORMAL_INIT_45_BIT_14_C : bit_vector(255 downto 0) := x"0A8E9A6A58F67B525ACAF0B7AD5BBF7E121B0A93A99097AAE7535B87A572FD6D";
   constant CPIX_NORMAL_INIT_46_BIT_00_C : bit_vector(255 downto 0) := x"26330906D7EC6DA7CC5B524F198ACC13659C70417F9AC993A4B5F2C2D7CA40F6";
   constant CPIX_NORMAL_INIT_46_BIT_01_C : bit_vector(255 downto 0) := x"8AFDA117E5E48DCE43A4D80C5C00BE427C36036990AF6B81B422EC3D4E3526F8";
   constant CPIX_NORMAL_INIT_46_BIT_02_C : bit_vector(255 downto 0) := x"CE36F3457EA4AA7E6CD617DDEC31EA8012A7EAEFAA0337016901ADA46F54C1C6";
   constant CPIX_NORMAL_INIT_46_BIT_03_C : bit_vector(255 downto 0) := x"03CEBFE2AD2A372C40E43C01EF05E8AA2C88B3E1D68D80DA4DD95E0DFB4D130A";
   constant CPIX_NORMAL_INIT_46_BIT_04_C : bit_vector(255 downto 0) := x"3BCF6F6BE65DE27903848533F3297D734503BAF7BC9BA65D9CDF7A15DA0015EF";
   constant CPIX_NORMAL_INIT_46_BIT_05_C : bit_vector(255 downto 0) := x"E12B6BE473047032F0777161012CC4D7A1FBD48273FE92008EE1C11331068FF3";
   constant CPIX_NORMAL_INIT_46_BIT_06_C : bit_vector(255 downto 0) := x"09C7942EA7785EA463018DA56261804995A4107FD294578FE901C1C89299DEFD";
   constant CPIX_NORMAL_INIT_46_BIT_07_C : bit_vector(255 downto 0) := x"508DE6459481E5769369A569A0C886C87E2716F50CBB72DF06E6E021F6F8EC2C";
   constant CPIX_NORMAL_INIT_46_BIT_08_C : bit_vector(255 downto 0) := x"084DDDCCEB882A31E120577423D6872EAAFCA4774DE33FF2EA4CC12052381A53";
   constant CPIX_NORMAL_INIT_46_BIT_09_C : bit_vector(255 downto 0) := x"148993FB1E8E3D90D829CDD5A6EE028555424DF52153417CAD42E6072FA18355";
   constant CPIX_NORMAL_INIT_46_BIT_10_C : bit_vector(255 downto 0) := x"A6CE9E7C1C7D49FA27D9164A0F5BF71AAB933AFFBE4A4A94D91809C9EF379540";
   constant CPIX_NORMAL_INIT_46_BIT_11_C : bit_vector(255 downto 0) := x"B85043B2F8D37875C5D7147FBC7DFF77665D83D7163C1F34DE5054BC2F5C42B2";
   constant CPIX_NORMAL_INIT_46_BIT_12_C : bit_vector(255 downto 0) := x"DBF8887D4A7B8B5DCC15B1A8DC55F97B1DD3EB4D57AA9DAAED39807D3DCCEDBD";
   constant CPIX_NORMAL_INIT_46_BIT_13_C : bit_vector(255 downto 0) := x"E3F13CF7ADB50045227D7BEB3715FB5AAA1C9AC811BE779A2BB6EE132DA21CC5";
   constant CPIX_NORMAL_INIT_46_BIT_14_C : bit_vector(255 downto 0) := x"0B6E00DE187F3EA0B533F14F653BF79A55F560CC1C7DCE15437B71AFA77ABCA7";
   constant CPIX_NORMAL_INIT_47_BIT_00_C : bit_vector(255 downto 0) := x"6B0D1F91859A78050FAEDA727FB5260680846EB28A705E4B74E0AC366697A7BB";
   constant CPIX_NORMAL_INIT_47_BIT_01_C : bit_vector(255 downto 0) := x"B3E15809315BDBB5CA135737E417BFC2D26FCEF750C34D36B18342B8EAB6927A";
   constant CPIX_NORMAL_INIT_47_BIT_02_C : bit_vector(255 downto 0) := x"4A7B474090FE48753B10716E5BA42B234855013E8515892CA2DCFD2B4ADFC982";
   constant CPIX_NORMAL_INIT_47_BIT_03_C : bit_vector(255 downto 0) := x"F98668B07AE699951C8DF8DA5D8043D0B93D03F96A038B927BC4565307B68578";
   constant CPIX_NORMAL_INIT_47_BIT_04_C : bit_vector(255 downto 0) := x"1B2272188528B9E47A77CCD8A353396EA81215357C23D46A920ED72E21B5F160";
   constant CPIX_NORMAL_INIT_47_BIT_05_C : bit_vector(255 downto 0) := x"670522F1D59E01C24B730B0714131D960B08003ECF2F144F986A7E7620249EFE";
   constant CPIX_NORMAL_INIT_47_BIT_06_C : bit_vector(255 downto 0) := x"0D67259C251D6FBEE3187FD30AC70D816D9E166F2C41F9EA753C512B60D63DE2";
   constant CPIX_NORMAL_INIT_47_BIT_07_C : bit_vector(255 downto 0) := x"6932C1B935FCCB012438083F25EC59FDB68FE4718E88B352EACB780B22A1C286";
   constant CPIX_NORMAL_INIT_47_BIT_08_C : bit_vector(255 downto 0) := x"E96AA8FDF951A5D8D69B65923EBA8839A7C7FD8CC25914A6D44433C6DA965831";
   constant CPIX_NORMAL_INIT_47_BIT_09_C : bit_vector(255 downto 0) := x"2D3CEF07FF3183009F28BFC8C5164401ADF72A9AAC2EE22B568AC8FEB90EE484";
   constant CPIX_NORMAL_INIT_47_BIT_10_C : bit_vector(255 downto 0) := x"1F0BF55793EAAC3FC5524C5FB9012021004E6E62B36A9B5A863984FD5F8D2E85";
   constant CPIX_NORMAL_INIT_47_BIT_11_C : bit_vector(255 downto 0) := x"151A2A2D22462E7C99745F2EC9F26AFD25F52020A9BA313535BF76817DED1D3B";
   constant CPIX_NORMAL_INIT_47_BIT_12_C : bit_vector(255 downto 0) := x"5033F2A654E47E7164306A54F5E246229FA9358EF955649388D811E63D26EBB1";
   constant CPIX_NORMAL_INIT_47_BIT_13_C : bit_vector(255 downto 0) := x"388ED46C82DD527B397576D573A615E1EBA665A52E1A0D505739A97B39B475CC";
   constant CPIX_NORMAL_INIT_47_BIT_14_C : bit_vector(255 downto 0) := x"44099981956F7B1B13DA9BBDAE48CB898D725295A5209182EE91B1705AE622C8";
   constant CPIX_NORMAL_INIT_48_BIT_00_C : bit_vector(255 downto 0) := x"96309D41606D37367086F6E42FE846432F962F8BAEAFBAEAB917CBD83371036D";
   constant CPIX_NORMAL_INIT_48_BIT_01_C : bit_vector(255 downto 0) := x"68F111BAC0C80C77F42B1E80FA9ABAFD3384DE3F7E74C3D03FB367606F0E85DC";
   constant CPIX_NORMAL_INIT_48_BIT_02_C : bit_vector(255 downto 0) := x"DBE5C09F3D156D4A2B6372F6CB82A325B5507DA1047CEB31B56936DBC71BA421";
   constant CPIX_NORMAL_INIT_48_BIT_03_C : bit_vector(255 downto 0) := x"9F29C0F54B69A1F618D88E50103D3236E0C36C776441DCD808A1EC77A3223F6B";
   constant CPIX_NORMAL_INIT_48_BIT_04_C : bit_vector(255 downto 0) := x"9340BAE56C63BA9144E1576CDDABB30A5F5632FF52A026692185186AE8D6FD46";
   constant CPIX_NORMAL_INIT_48_BIT_05_C : bit_vector(255 downto 0) := x"5E1B9FB6144604867DA89E3CAFCC554A51C54184D57B595D8AB65FA49502D571";
   constant CPIX_NORMAL_INIT_48_BIT_06_C : bit_vector(255 downto 0) := x"ED2678467B30D703FDA7CF5715B28B73D47175ABA1F730AA1BD0F2898ADF2F7B";
   constant CPIX_NORMAL_INIT_48_BIT_07_C : bit_vector(255 downto 0) := x"0C9DE8017B22F9CB18299A25F4C828981E637BDBA04CED7CDF64BF371CEA2243";
   constant CPIX_NORMAL_INIT_48_BIT_08_C : bit_vector(255 downto 0) := x"12A8F3D470377A4026957B9A29A56DD3A5E9055AB701CF1D1627EB63E4A70F2D";
   constant CPIX_NORMAL_INIT_48_BIT_09_C : bit_vector(255 downto 0) := x"F8AECC978E3DB1B909B5A9F77976EEE5612D2E7C1568EFC0320355B403CED46F";
   constant CPIX_NORMAL_INIT_48_BIT_10_C : bit_vector(255 downto 0) := x"B3B060BFFCAA190E9173CF7D497FFE5704BC92A55D3AEF47C5DF8350DC3650BE";
   constant CPIX_NORMAL_INIT_48_BIT_11_C : bit_vector(255 downto 0) := x"9771C1EE01FFDFBCFF88304332872CD6EA965D1C939BFD044F788542195D9B8F";
   constant CPIX_NORMAL_INIT_48_BIT_12_C : bit_vector(255 downto 0) := x"1E9AB61C11CC9A9FAFE1FB915F0DDD59375A27453A95CD873B12367F66ACCC5D";
   constant CPIX_NORMAL_INIT_48_BIT_13_C : bit_vector(255 downto 0) := x"74767A873D4C466B91E8440EF094E807EBC3343E6B495D6AF139B2B49E9FD817";
   constant CPIX_NORMAL_INIT_48_BIT_14_C : bit_vector(255 downto 0) := x"8C189884569ADF1B441B029BD71D6367AF69D1A9B337614915168CDE3336B692";
   constant CPIX_NORMAL_INIT_49_BIT_00_C : bit_vector(255 downto 0) := x"0D95D3C3A3EA49C3CECC2E39C0853214C2C551D5AB3A606E3F1AAE5A588513BE";
   constant CPIX_NORMAL_INIT_49_BIT_01_C : bit_vector(255 downto 0) := x"81FE7515515A0AEA92A5A64CCFFB14EA3A718CC1E357DBE6B09F74DCA4DB90EE";
   constant CPIX_NORMAL_INIT_49_BIT_02_C : bit_vector(255 downto 0) := x"8866EDF2806557BC58A393211F3E1582BD5E0692F86B5BEAD8911EF9A2CE3F54";
   constant CPIX_NORMAL_INIT_49_BIT_03_C : bit_vector(255 downto 0) := x"2F0EADBD6A1B78732159F48ADD3A3FA7ED13AC582DF2797168BAB6F931EB2966";
   constant CPIX_NORMAL_INIT_49_BIT_04_C : bit_vector(255 downto 0) := x"0C1E3F4941899A7FFC1AFF0C647D51106B5E1D2EDF227F40E92C6CB83872D303";
   constant CPIX_NORMAL_INIT_49_BIT_05_C : bit_vector(255 downto 0) := x"DEB165F9102CC95ABA3351AD399772AC851A4EEDD8D08047AC15B5649FFC587A";
   constant CPIX_NORMAL_INIT_49_BIT_06_C : bit_vector(255 downto 0) := x"060E029C34D9B0C6B42A9DDB2430742C44F1C65B497C30A9D1ABA003D2B8A406";
   constant CPIX_NORMAL_INIT_49_BIT_07_C : bit_vector(255 downto 0) := x"05129F51F028EB4F15DC2AC99493A11161A3DCA896301FB0A1C82A02C01887F8";
   constant CPIX_NORMAL_INIT_49_BIT_08_C : bit_vector(255 downto 0) := x"F5D55C3859B55F3860EEAAA53B0D355E8F9D2F84E365EF52E657F6FD14C6ABCF";
   constant CPIX_NORMAL_INIT_49_BIT_09_C : bit_vector(255 downto 0) := x"6F07494B8EE5AD3AED5B84156DC744E28DAC913EAFF6D357CEBEDDFD7C577A37";
   constant CPIX_NORMAL_INIT_49_BIT_10_C : bit_vector(255 downto 0) := x"5C959F203DC27DF8415CC2D8E9864AED8D813D7A7A8DC7ACEA45A7751937DBCD";
   constant CPIX_NORMAL_INIT_49_BIT_11_C : bit_vector(255 downto 0) := x"5247D2B5CC59D960737CDD0E7344B0B4F7CEACB352AEA7CD5875E77D978773A5";
   constant CPIX_NORMAL_INIT_49_BIT_12_C : bit_vector(255 downto 0) := x"7B9428E37A714D445045504EAD957A88CCA6EBA28C75A77A435CCE7FB58EB73F";
   constant CPIX_NORMAL_INIT_49_BIT_13_C : bit_vector(255 downto 0) := x"4C3D8954A3C3BDA3B74A3F1E4A856259D5768542ACAC33C3D2B4EC7DDE35321D";
   constant CPIX_NORMAL_INIT_49_BIT_14_C : bit_vector(255 downto 0) := x"030D7CE7138A3C4578D20BF97AFCD98644E9E729CCCEA3A27305AC779A8D84F6";
   constant CPIX_NORMAL_INIT_4A_BIT_00_C : bit_vector(255 downto 0) := x"3AE5CAFE89EF33E07E3CA8237AC7D2241C28139E84B436347E3B836FA0832315";
   constant CPIX_NORMAL_INIT_4A_BIT_01_C : bit_vector(255 downto 0) := x"97185E8F29E41E8F173A6316E938BF69B3F613EBC08DB2B30AF74C96F817BFCE";
   constant CPIX_NORMAL_INIT_4A_BIT_02_C : bit_vector(255 downto 0) := x"89CBD20E01F0FE0EA0EA6337B1BD63C1CCF20418534838934A6BE9A3F3D6C1AA";
   constant CPIX_NORMAL_INIT_4A_BIT_03_C : bit_vector(255 downto 0) := x"5D2C93394B474B177CD2521C953A81E72ABBDCC95018AFF217B2B89CFD739C2F";
   constant CPIX_NORMAL_INIT_4A_BIT_04_C : bit_vector(255 downto 0) := x"45DED78DF1858F9E31544B1283EABA3A639A5F20F2E697835983BDD36A320220";
   constant CPIX_NORMAL_INIT_4A_BIT_05_C : bit_vector(255 downto 0) := x"9C35515DA8A1E9A0EE74747D33D23FA38D0C1966E4D9E01D70A1300990A53D3F";
   constant CPIX_NORMAL_INIT_4A_BIT_06_C : bit_vector(255 downto 0) := x"0A57C88361A188C4823686EEEC4DEB91EB08AED698102079F726D4589C90881F";
   constant CPIX_NORMAL_INIT_4A_BIT_07_C : bit_vector(255 downto 0) := x"76C2C3FC9D6F54CB31E9AE84514BF398D9B162863597D54ED460F50E8051F993";
   constant CPIX_NORMAL_INIT_4A_BIT_08_C : bit_vector(255 downto 0) := x"BD5E4CE883F3F6E680EFFDD1D2FD09DE4F479C080D375DBF6AB679357A8927F2";
   constant CPIX_NORMAL_INIT_4A_BIT_09_C : bit_vector(255 downto 0) := x"8DC0F4216D2C3686ED1DD45D716E371ABE354A57C310CE66E0EDE2D491B62C46";
   constant CPIX_NORMAL_INIT_4A_BIT_10_C : bit_vector(255 downto 0) := x"DA149EAD06BA25919C2BC2D32FE6D98C071CE0431055CF66845336D255849B23";
   constant CPIX_NORMAL_INIT_4A_BIT_11_C : bit_vector(255 downto 0) := x"90C6DBC5B3599C0265FB75891CA66FB24EEBE5AAB8BC67CF259CC09854E45A56";
   constant CPIX_NORMAL_INIT_4A_BIT_12_C : bit_vector(255 downto 0) := x"0ED2B83AA5CD13D3D2A56C9E52871A6E2FF2BC29E2464D3C0B7DAF3CAFEA84EA";
   constant CPIX_NORMAL_INIT_4A_BIT_13_C : bit_vector(255 downto 0) := x"64B96C4AEE8D1B6BED82B5906644FB8033E37D06037BEC041F34E3CAEBCB47F4";
   constant CPIX_NORMAL_INIT_4A_BIT_14_C : bit_vector(255 downto 0) := x"2524932855C4F2B0C55D293126FEBE7B64E3267183A33C5CF6325773AB327D72";
   constant CPIX_NORMAL_INIT_4B_BIT_00_C : bit_vector(255 downto 0) := x"2AAAE496DC6D1144412BDD9C7562D7086F029F88CCBC5C7832935DA297925723";
   constant CPIX_NORMAL_INIT_4B_BIT_01_C : bit_vector(255 downto 0) := x"B1AA62E9A99DBF75C224686005D1562CA3DBFE3128A0BDB20FD6EE0A0DF3666C";
   constant CPIX_NORMAL_INIT_4B_BIT_02_C : bit_vector(255 downto 0) := x"333C829A130D660DA5E057435E09CCBD0C97DBFF47C8750E78BC10806024ECAD";
   constant CPIX_NORMAL_INIT_4B_BIT_03_C : bit_vector(255 downto 0) := x"89A5CB94995E2A3E4215B2EB100746D64D4366E92EF3A018C425137BD5F8CB42";
   constant CPIX_NORMAL_INIT_4B_BIT_04_C : bit_vector(255 downto 0) := x"766DC9A278611E1793877953F50C86890A40301EC40B604D7BC9253727C7CE79";
   constant CPIX_NORMAL_INIT_4B_BIT_05_C : bit_vector(255 downto 0) := x"1E722789E5B57A15A208F373467A0F9A4825C8AB6D52C52004667449E6C7B22F";
   constant CPIX_NORMAL_INIT_4B_BIT_06_C : bit_vector(255 downto 0) := x"682E337BA3FC69EA4EEDDC406239534E9C359378E06B1C38E9DD300754ABD44C";
   constant CPIX_NORMAL_INIT_4B_BIT_07_C : bit_vector(255 downto 0) := x"0B0E5E2811204274EEB88564F258ED7D649EE8A62EB17BDADCD31E490622CBAB";
   constant CPIX_NORMAL_INIT_4B_BIT_08_C : bit_vector(255 downto 0) := x"1C5BC849D68D34C61ED388454F4608DC09B827CBFCE06F7507784A19523C3BEB";
   constant CPIX_NORMAL_INIT_4B_BIT_09_C : bit_vector(255 downto 0) := x"470B41D2CD46410EDD1A6E22EF24CAB817190A7D710D5A74F03885757E857F3B";
   constant CPIX_NORMAL_INIT_4B_BIT_10_C : bit_vector(255 downto 0) := x"EF62A07B6C679A542C00623B30CAFBDCAA10FE5FA6DFF8FDE857FCDFA76A9410";
   constant CPIX_NORMAL_INIT_4B_BIT_11_C : bit_vector(255 downto 0) := x"C4541DCEE1E70E0E7ECC59C97CFCBD003EC387297CD678D23490B43EE8124EFE";
   constant CPIX_NORMAL_INIT_4B_BIT_12_C : bit_vector(255 downto 0) := x"A5F5D1191626B9C2F7C3DF3B62BD3E3B3CC7C6A0841AEE94EFD9A7105A21E441";
   constant CPIX_NORMAL_INIT_4B_BIT_13_C : bit_vector(255 downto 0) := x"85BC82FEEADE4A6700CE446E339E64FB47A118AB1BD5C8FF192DD381638237A0";
   constant CPIX_NORMAL_INIT_4B_BIT_14_C : bit_vector(255 downto 0) := x"62A653AA6A1542AAF56C54ABE7CBB0166CEDEE38AA4DAC54A8CA57AB9DDA9B94";
   constant CPIX_NORMAL_INIT_4C_BIT_00_C : bit_vector(255 downto 0) := x"59822E1CC69C0F8DAA35FDBC2431B6330E6DB00907C6F0963424BE23945B052E";
   constant CPIX_NORMAL_INIT_4C_BIT_01_C : bit_vector(255 downto 0) := x"F675DC455B539978DD732BD89B91D96C94D7A8EFD7B883B7AA6B5A0A835A8B97";
   constant CPIX_NORMAL_INIT_4C_BIT_02_C : bit_vector(255 downto 0) := x"66E40A87B199632276B4D17201CB728648AB4D3B41890F372BA59E77244F33E8";
   constant CPIX_NORMAL_INIT_4C_BIT_03_C : bit_vector(255 downto 0) := x"0D05CA65896305C1E2DA12E952F481C92868347B2CBB34DE320B2558593E1B3F";
   constant CPIX_NORMAL_INIT_4C_BIT_04_C : bit_vector(255 downto 0) := x"42C7D7C34F8212758295130312AE6EF4B15F537A197CE0EC6F48F86E920316F1";
   constant CPIX_NORMAL_INIT_4C_BIT_05_C : bit_vector(255 downto 0) := x"9AAACC16DDA5A187A449AD4BEDC74CAD4867DE93E8124F88AC8165E016BCF8F2";
   constant CPIX_NORMAL_INIT_4C_BIT_06_C : bit_vector(255 downto 0) := x"F8F8EDD93BFEBB32FAF22C180B3AAB71905D76D34324EB3051182DD335FE68D3";
   constant CPIX_NORMAL_INIT_4C_BIT_07_C : bit_vector(255 downto 0) := x"3FB0B1F64A3DFA7B7D63688820F12C9EEF421CFD58FB313670E043877B7238B6";
   constant CPIX_NORMAL_INIT_4C_BIT_08_C : bit_vector(255 downto 0) := x"5B28DE74C43BEE5C00BB7A3D7C24A28FC3111DE6624C3AE7213678FE255D645A";
   constant CPIX_NORMAL_INIT_4C_BIT_09_C : bit_vector(255 downto 0) := x"5AAD7E9B3CAFA39E075D629A31EDBFE5A8B44A5248CD33734FAD1FE95321771B";
   constant CPIX_NORMAL_INIT_4C_BIT_10_C : bit_vector(255 downto 0) := x"778E6450FE692196E4126A115156EEE3316C7042570B2CF976D66D733C36719F";
   constant CPIX_NORMAL_INIT_4C_BIT_11_C : bit_vector(255 downto 0) := x"3905FFC4683126D722450BE2596DF0085FFB57352A517832F5C3A7A4CAE5B223";
   constant CPIX_NORMAL_INIT_4C_BIT_12_C : bit_vector(255 downto 0) := x"64520C707DEE6254A74249DF60F50806FB87E53DC4C8B6A37C815870D5CBF393";
   constant CPIX_NORMAL_INIT_4C_BIT_13_C : bit_vector(255 downto 0) := x"7384A208DD2B2659D5D990A990AE985C5BCEEC2A0251DD2B0BB7CB1E4E9A9AEE";
   constant CPIX_NORMAL_INIT_4C_BIT_14_C : bit_vector(255 downto 0) := x"598EECA504AB65C0DCC4D7EF46D501E224A6BAAF6513AA4E6D52D24A09848748";
   constant CPIX_NORMAL_INIT_4D_BIT_00_C : bit_vector(255 downto 0) := x"737835AE2802CB45FA024D3E9AE044DC176DE3D54A51E12E873D3221F2972C13";
   constant CPIX_NORMAL_INIT_4D_BIT_01_C : bit_vector(255 downto 0) := x"A609867A6249F477A771FA5FCA7476E0C94644F7089E06FC3F802A092EF17E30";
   constant CPIX_NORMAL_INIT_4D_BIT_02_C : bit_vector(255 downto 0) := x"1440D9B17AC79F19E1FC91E054A4A689A1D80F242E35F2DF2357D8BD642FA040";
   constant CPIX_NORMAL_INIT_4D_BIT_03_C : bit_vector(255 downto 0) := x"D0DCC51FD4BBEBBFC465164F3412A00111A6BDFD53B5462B2D204D597EBBE795";
   constant CPIX_NORMAL_INIT_4D_BIT_04_C : bit_vector(255 downto 0) := x"CF258CBE4DDF93C303BACA64AE3AF4071937ED17440ECEC5D0D249483475936A";
   constant CPIX_NORMAL_INIT_4D_BIT_05_C : bit_vector(255 downto 0) := x"BD38C6BD7719E67849292E7468936E4D57A44956FBEBA39787C3AE7AE68483AD";
   constant CPIX_NORMAL_INIT_4D_BIT_06_C : bit_vector(255 downto 0) := x"77C36D15116FC83B03AAD591B433AF834F28D3A47CF44BAC466DCBF7BFE38445";
   constant CPIX_NORMAL_INIT_4D_BIT_07_C : bit_vector(255 downto 0) := x"E81A1A77685611C66E2DC3865D7F22607B935E809571FE70C5EF6B70A70A0A37";
   constant CPIX_NORMAL_INIT_4D_BIT_08_C : bit_vector(255 downto 0) := x"AB66B7A20211D0899E85FEF81E5F479AA6C98F1247F325FA0EE91688D16EC0EF";
   constant CPIX_NORMAL_INIT_4D_BIT_09_C : bit_vector(255 downto 0) := x"555D16D88DFC79B5CB6590FE17809E15743833D1B3FFF84B59B0033CC23FA07F";
   constant CPIX_NORMAL_INIT_4D_BIT_10_C : bit_vector(255 downto 0) := x"396FC12302699BEFD1FD31F726BF220BA795A0A809F0DE123F752A170D531A33";
   constant CPIX_NORMAL_INIT_4D_BIT_11_C : bit_vector(255 downto 0) := x"39C67767E8EB07DF81F75D0D5704C0489E1692DF9E645134631A7A8B6F16BF73";
   constant CPIX_NORMAL_INIT_4D_BIT_12_C : bit_vector(255 downto 0) := x"A0DE2BFE1BB3F868083C63F038D789E7C977F1E653788391CAF460E22CB7F410";
   constant CPIX_NORMAL_INIT_4D_BIT_13_C : bit_vector(255 downto 0) := x"0DFB2C6E33CD47FDF9259922A559B731F3506D1D4C369D04E373E215BE3447B8";
   constant CPIX_NORMAL_INIT_4D_BIT_14_C : bit_vector(255 downto 0) := x"B8861C570E1A2A52B686F1B4535A8618517A8A5A96F85D5F0EF6954F0FF9106E";
   constant CPIX_NORMAL_INIT_4E_BIT_00_C : bit_vector(255 downto 0) := x"428DD1D7352D33CAF3337A34083D415785D09E1DD15F9D71112BBDF6F71CBB8B";
   constant CPIX_NORMAL_INIT_4E_BIT_01_C : bit_vector(255 downto 0) := x"C1F371E2AC445324EBF5A2E1FEC41F54B4CABDE6BF8CD109CD5D293612C584F1";
   constant CPIX_NORMAL_INIT_4E_BIT_02_C : bit_vector(255 downto 0) := x"91F55EE70A63EC6644431BB7EECD4EFE72C2A97577B5E9B2A9AC828F22158F4D";
   constant CPIX_NORMAL_INIT_4E_BIT_03_C : bit_vector(255 downto 0) := x"5FA506E96DC31708F3CC6EDDE401AC1F12F2F7F436F2249C4D1FB004F42A279C";
   constant CPIX_NORMAL_INIT_4E_BIT_04_C : bit_vector(255 downto 0) := x"59A732E8E21AD0358CA28BAA379A52BC85EF1B66D7CACE5379977237CDB66CD6";
   constant CPIX_NORMAL_INIT_4E_BIT_05_C : bit_vector(255 downto 0) := x"4BA2B33DF908F0C8C97866E1E4FF63401ECE2BD94ED949B63A8465EF67B9F478";
   constant CPIX_NORMAL_INIT_4E_BIT_06_C : bit_vector(255 downto 0) := x"33286E2EF0E74043C535EA3F6CD9C0AF4F61D7B7625920A17D654A40CB0F5EE8";
   constant CPIX_NORMAL_INIT_4E_BIT_07_C : bit_vector(255 downto 0) := x"452C9D17E9A20AB1DBD06D5AA45343399CAE8E799D21EEFE7A05AAE934FD258D";
   constant CPIX_NORMAL_INIT_4E_BIT_08_C : bit_vector(255 downto 0) := x"92E77AE5D69873A71DF9F4F48B36620D4A8D28EEB7BEED7791C147A5C4824988";
   constant CPIX_NORMAL_INIT_4E_BIT_09_C : bit_vector(255 downto 0) := x"648BC268763D262B14774DFBC92589D48432549A3D0DC3BCAA686EC7963087A3";
   constant CPIX_NORMAL_INIT_4E_BIT_10_C : bit_vector(255 downto 0) := x"C1983C2F04765ADD5486123BB85025CBD3C547365E95D9746DCEF41CB510E849";
   constant CPIX_NORMAL_INIT_4E_BIT_11_C : bit_vector(255 downto 0) := x"3F2F03B3056C3362807C496E0CEAF07D842423A4F5D1685DF15447E9DBD071C2";
   constant CPIX_NORMAL_INIT_4E_BIT_12_C : bit_vector(255 downto 0) := x"48CF77858F13A54A78AD07BE018B6385F304D0B274BEDA7561DDA35152CFF0D0";
   constant CPIX_NORMAL_INIT_4E_BIT_13_C : bit_vector(255 downto 0) := x"14B34F5953AB9D8E9FD40349CA69AE473FDAAC1F4CDCE29506BB4DDA6A1B079E";
   constant CPIX_NORMAL_INIT_4E_BIT_14_C : bit_vector(255 downto 0) := x"53236BB7FA7A2D1F6CFAB939FFD0FC025AFACC8C0D35F2C2F045DBE2F185E3FF";
   constant CPIX_NORMAL_INIT_4F_BIT_00_C : bit_vector(255 downto 0) := x"4E16253701184FA3CBFFDD496C482C6B50FB6C1A7DCFC048205A3FD6DF2E5151";
   constant CPIX_NORMAL_INIT_4F_BIT_01_C : bit_vector(255 downto 0) := x"9AB4D5E4513AD66EAF1B4B3CBBFFEA0AE8DDE3B7D5EAD1F598C905A3C503F96D";
   constant CPIX_NORMAL_INIT_4F_BIT_02_C : bit_vector(255 downto 0) := x"602B2001B91F02E57C2A514D5F184074B9C17A445E99C62341F8D748E26D3BE6";
   constant CPIX_NORMAL_INIT_4F_BIT_03_C : bit_vector(255 downto 0) := x"F7D94D3BABEFFF9690A7CF402F60632982BC223876631B83434FE7DB359F06BC";
   constant CPIX_NORMAL_INIT_4F_BIT_04_C : bit_vector(255 downto 0) := x"5A1818FB4B14B1C342C8736E4678880B1C6A03753F53CC5346C5D94C373B796C";
   constant CPIX_NORMAL_INIT_4F_BIT_05_C : bit_vector(255 downto 0) := x"ED6C23D54B9D06394C73F45580E61CC419ADD912C3A12B5BA73C5E3CA728E386";
   constant CPIX_NORMAL_INIT_4F_BIT_06_C : bit_vector(255 downto 0) := x"613BE1E115670D79602A03136CDF365AABE05D7B08662C6E5C39D99F768D3B19";
   constant CPIX_NORMAL_INIT_4F_BIT_07_C : bit_vector(255 downto 0) := x"61494B880A3FE3ADF97830FE18F33FA9D670FB9FBC2DFE255906624DDB8B4356";
   constant CPIX_NORMAL_INIT_4F_BIT_08_C : bit_vector(255 downto 0) := x"6E17E62F08044BBF7F2F308568ED122582CEA90745AC41037B20ED9D5EC15393";
   constant CPIX_NORMAL_INIT_4F_BIT_09_C : bit_vector(255 downto 0) := x"4356CD29D5CE26A669B0518A083EF70E49ED91425523E90C90EE51E90DD2E6A6";
   constant CPIX_NORMAL_INIT_4F_BIT_10_C : bit_vector(255 downto 0) := x"135CBA778F6608E31DC830B6106F487D1722F00F759FD7DC32602DE090B0F941";
   constant CPIX_NORMAL_INIT_4F_BIT_11_C : bit_vector(255 downto 0) := x"4B9E9A9CF16865B921FE6010415D0676AE0641553892EF433781E73E7886D2EE";
   constant CPIX_NORMAL_INIT_4F_BIT_12_C : bit_vector(255 downto 0) := x"401D0C7CBE321E9F649109A610D63A0180516773274B61F047DF4D5BC369ADC6";
   constant CPIX_NORMAL_INIT_4F_BIT_13_C : bit_vector(255 downto 0) := x"490E60F0747C023A334A3FD64F75597495F1688B465108550A85F9E5DB4F0B03";
   constant CPIX_NORMAL_INIT_4F_BIT_14_C : bit_vector(255 downto 0) := x"09419068794B2FADA8E3D14ABF05E8E5C07E5C050D462152153D5EF810AC2456";
   constant CPIX_NORMAL_INIT_50_BIT_00_C : bit_vector(255 downto 0) := x"8054F9CE7EF765854A25FC6C971DC10B1F9D69871F15E2EB878417DA7E2147FA";
   constant CPIX_NORMAL_INIT_50_BIT_01_C : bit_vector(255 downto 0) := x"17004439B9A627BC63A696FBA62236C732DF95D901B885E4CA080C589B1E3BC2";
   constant CPIX_NORMAL_INIT_50_BIT_02_C : bit_vector(255 downto 0) := x"F889D0E396D1FE6680EFA0B3EA307B75F135755CF76FADE9C03D95756AE7E8FF";
   constant CPIX_NORMAL_INIT_50_BIT_03_C : bit_vector(255 downto 0) := x"E1CADA609D4D189F565D3C717BFF52F77BB0A2BD450683A40DC8C523504C9AEF";
   constant CPIX_NORMAL_INIT_50_BIT_04_C : bit_vector(255 downto 0) := x"7E9BA98E0C31B720A293FE81017231E38791436B8271C6C118615F92C66BB75B";
   constant CPIX_NORMAL_INIT_50_BIT_05_C : bit_vector(255 downto 0) := x"661EB7DE7BC3F8C2F6CA44047A3D3C268BEB0CCCE535EA95BAE1D537CE05F535";
   constant CPIX_NORMAL_INIT_50_BIT_06_C : bit_vector(255 downto 0) := x"65CA8B9FBCDFA098B780D9FD31D803184E50E8A3960048114BC1BAFC95D5FFE5";
   constant CPIX_NORMAL_INIT_50_BIT_07_C : bit_vector(255 downto 0) := x"CEFBA190E10370D1AAADDA1660E0D9DE14CC3FC5F4EB927D3ECA40E650A98CFF";
   constant CPIX_NORMAL_INIT_50_BIT_08_C : bit_vector(255 downto 0) := x"DB3D572E765915120FC020C27D024357BBF0BD6B41BDEDCDEC36E52DC1EB9CFB";
   constant CPIX_NORMAL_INIT_50_BIT_09_C : bit_vector(255 downto 0) := x"C673A8CD98B90ADDF601D64EC1CFCD02EB9885B856753A33F27D5161DB34B6E9";
   constant CPIX_NORMAL_INIT_50_BIT_10_C : bit_vector(255 downto 0) := x"5187498EE8C6587C2CB0D299D3AF200087022BC6147805FDA88A7ED9A263DCE5";
   constant CPIX_NORMAL_INIT_50_BIT_11_C : bit_vector(255 downto 0) := x"526E011D312CA8E867FF7DF07A74BB29A04E0AE74CEAFCA2595623DD18EDAC31";
   constant CPIX_NORMAL_INIT_50_BIT_12_C : bit_vector(255 downto 0) := x"FFA8DE79472527FF374DB5BB354BF4C0464873DA5A0CD92A674E65CAAC19EC53";
   constant CPIX_NORMAL_INIT_50_BIT_13_C : bit_vector(255 downto 0) := x"9D4DD76A06036CDC745DC27A84BB6477302FE21A736EDE3E8CB63C16B3CE0AD9";
   constant CPIX_NORMAL_INIT_50_BIT_14_C : bit_vector(255 downto 0) := x"C75AF643B551456D395B855CB01AA5DB7997A7E48DF4409CF3FE3DEFA0301553";
   constant CPIX_NORMAL_INIT_51_BIT_00_C : bit_vector(255 downto 0) := x"5F694AF00229823734C539C369E738C2D32CCD4E545EC9637EC0A8A72163A32B";
   constant CPIX_NORMAL_INIT_51_BIT_01_C : bit_vector(255 downto 0) := x"2600C0C36C692DD5C8BBB7775A6A7CCD48E3DD34B02199284A136A00A2058570";
   constant CPIX_NORMAL_INIT_51_BIT_02_C : bit_vector(255 downto 0) := x"12A32C065A1D00E1E5399847CB7728A9E339E523CB8C056868DD91C7D454A0DA";
   constant CPIX_NORMAL_INIT_51_BIT_03_C : bit_vector(255 downto 0) := x"C08F9AC4BF1FCBA78C75991747F0515502A7441F2883602D6AD1AD7CA494DE9D";
   constant CPIX_NORMAL_INIT_51_BIT_04_C : bit_vector(255 downto 0) := x"CA4CB27C27918CFD5502D7D819D3BB8C4819CFB5C855A8AFD96E99E75BEBB78D";
   constant CPIX_NORMAL_INIT_51_BIT_05_C : bit_vector(255 downto 0) := x"53E475BE42588A8B54CA2D4378A817C7C672E506566BE340258189F3B5915BA4";
   constant CPIX_NORMAL_INIT_51_BIT_06_C : bit_vector(255 downto 0) := x"56766F15691CEDAD58685511CBAD54BB95241127FBBE5001E91553C5352AD1A1";
   constant CPIX_NORMAL_INIT_51_BIT_07_C : bit_vector(255 downto 0) := x"67E5234F930E19919196D5009B3B01A05F0E440FC3DCB01F12E8EBDB6E3F5F4B";
   constant CPIX_NORMAL_INIT_51_BIT_08_C : bit_vector(255 downto 0) := x"43F6B6A35C388C2A1C434E64235E04ABC99605776C333007023BFC3C837EB39D";
   constant CPIX_NORMAL_INIT_51_BIT_09_C : bit_vector(255 downto 0) := x"65F4CC61720182C09F8E9701C7764157C7565E1A982395E904362367032E5922";
   constant CPIX_NORMAL_INIT_51_BIT_10_C : bit_vector(255 downto 0) := x"DFC363D100CE33D10AB6787E7B82E57CA0C1D5F5F2466EFBFF86E2D629BBBDF8";
   constant CPIX_NORMAL_INIT_51_BIT_11_C : bit_vector(255 downto 0) := x"E102EC63706FF9DFA6BB7BBF37AEAA62EF07F342191863F87FD833A4CC73335A";
   constant CPIX_NORMAL_INIT_51_BIT_12_C : bit_vector(255 downto 0) := x"B88B22C0DCF32CC7E3373CBFF5CC73C796B8271196AC96FD3BC89DA58CB7A8E0";
   constant CPIX_NORMAL_INIT_51_BIT_13_C : bit_vector(255 downto 0) := x"883BFBCD4526F7EC7B713DFE28EE63491D1D7DCA63238CED648DE96AFD832788";
   constant CPIX_NORMAL_INIT_51_BIT_14_C : bit_vector(255 downto 0) := x"1DDFEF056B4C3E8042B8FD7EF0B37D6908AE8B7EB36C7D6D73BF279610D2F626";
   constant CPIX_NORMAL_INIT_52_BIT_00_C : bit_vector(255 downto 0) := x"029C5ECC4C2ABCED925CA1988E2AB5177D45031A1F60E29EAD1E88416518F6F5";
   constant CPIX_NORMAL_INIT_52_BIT_01_C : bit_vector(255 downto 0) := x"3E80FF8784F19F8F16B6199212E4CD43901F6F874E8345C7C1FC675434590BB9";
   constant CPIX_NORMAL_INIT_52_BIT_02_C : bit_vector(255 downto 0) := x"DC51B214BBBD378E4EDE1E67302FD8A79601F26BAC1FFEC912083D11D97ED0C8";
   constant CPIX_NORMAL_INIT_52_BIT_03_C : bit_vector(255 downto 0) := x"4AE28B96D183086AC9C1B2E7298222FAD73A1AEE7E6C6F15D35E87AA034213C5";
   constant CPIX_NORMAL_INIT_52_BIT_04_C : bit_vector(255 downto 0) := x"9C9B5DC58A90D7596D56F6486C8DDF22BD5BAE3C60CC06ACC91319DCEBC158AC";
   constant CPIX_NORMAL_INIT_52_BIT_05_C : bit_vector(255 downto 0) := x"AD7B0F2291E40911BF143BED4C33999D2786BFF861A138EABE80CB4CD4BF2C4F";
   constant CPIX_NORMAL_INIT_52_BIT_06_C : bit_vector(255 downto 0) := x"0764183C3E9A79983150301742A3CAA302B88D283369D1A048EDD6E7BD78E937";
   constant CPIX_NORMAL_INIT_52_BIT_07_C : bit_vector(255 downto 0) := x"48C224A720BEB90586D9C0DEF0FC8C3F6F85E1B758AE402631CD99829F06CF81";
   constant CPIX_NORMAL_INIT_52_BIT_08_C : bit_vector(255 downto 0) := x"B198B142650763ADE0781FB6587F2F96FAFE01DE74563B858EB83E5756D79515";
   constant CPIX_NORMAL_INIT_52_BIT_09_C : bit_vector(255 downto 0) := x"5644E042F3DAA79F49487BCEB36012E0551673504E6F2FBB833F77E152C49E49";
   constant CPIX_NORMAL_INIT_52_BIT_10_C : bit_vector(255 downto 0) := x"431A038E2B3B3B4AA927934C61B43ACDBCCE62415E9417FDE38CF77B29E576AA";
   constant CPIX_NORMAL_INIT_52_BIT_11_C : bit_vector(255 downto 0) := x"2C508DAC95AAAA228DF87D8614A5628A9B3CECCAC385B7DDF47EC9922EFC64FD";
   constant CPIX_NORMAL_INIT_52_BIT_12_C : bit_vector(255 downto 0) := x"7F8CDF3B902276912A5F929869067640E1B49878043663CFAACB5FDFE5B5EB03";
   constant CPIX_NORMAL_INIT_52_BIT_13_C : bit_vector(255 downto 0) := x"622100E359F3DD4C301D4E0CDC70E456365DCE13E40DA3BBA9C1C0A15A5CFABB";
   constant CPIX_NORMAL_INIT_52_BIT_14_C : bit_vector(255 downto 0) := x"0C30C95A12120DEE4CCA772B135AAF6E59C9A7AC1504D39228AF33F55DF5E2EA";
   constant CPIX_NORMAL_INIT_53_BIT_00_C : bit_vector(255 downto 0) := x"27657D01B2D02ECF1FDCFA376BFFDEEDEC058682D73479B3C2253E3B194A89B4";
   constant CPIX_NORMAL_INIT_53_BIT_01_C : bit_vector(255 downto 0) := x"5317890FC8306AA283F38E717332896CEDE484D7BCDD3EC5460109034E18E798";
   constant CPIX_NORMAL_INIT_53_BIT_02_C : bit_vector(255 downto 0) := x"42E604ED108106BE7AE39163F4C4C859627BE856D8E645D547F5A75B594FBC84";
   constant CPIX_NORMAL_INIT_53_BIT_03_C : bit_vector(255 downto 0) := x"B5589448229D5550D3BF4372DEA2F0CEC7D799F757354372175428A64332326F";
   constant CPIX_NORMAL_INIT_53_BIT_04_C : bit_vector(255 downto 0) := x"AB6D0C2987F31CFCDA88048A0CC37B2A123DE07FE705A4FC1B4B3D80BEE0689B";
   constant CPIX_NORMAL_INIT_53_BIT_05_C : bit_vector(255 downto 0) := x"47733B00DE576A444D48613487368572E3F2D267C6D3524580D515511B2434AA";
   constant CPIX_NORMAL_INIT_53_BIT_06_C : bit_vector(255 downto 0) := x"75D7073A4F00BF9FC09173315F31D058D7D3CFF34CA41791A7EEA267BB46C7E3";
   constant CPIX_NORMAL_INIT_53_BIT_07_C : bit_vector(255 downto 0) := x"5435EABDAF99C1D64F43E63783D291B52B2C94B2F8FA5643EE3BD0324BBE85EA";
   constant CPIX_NORMAL_INIT_53_BIT_08_C : bit_vector(255 downto 0) := x"3107D9190545C79F99ADFA6110E7D5044C391AB4167618C1CA323B817C096A72";
   constant CPIX_NORMAL_INIT_53_BIT_09_C : bit_vector(255 downto 0) := x"65C06C2C5CD48D6010B1B7562AD601A5FA6F5ACBAFF9E6339B9672DD221F5DDF";
   constant CPIX_NORMAL_INIT_53_BIT_10_C : bit_vector(255 downto 0) := x"EB41CA93C9FE84AD692B8BA5D6BE4AE1D51DFF31706AF37BC29623E1C8D3A7AF";
   constant CPIX_NORMAL_INIT_53_BIT_11_C : bit_vector(255 downto 0) := x"6AC7627207A5D688D74C240B04F3E5ECCD177DC0AB8E696FDC3314D8FF3AD419";
   constant CPIX_NORMAL_INIT_53_BIT_12_C : bit_vector(255 downto 0) := x"32AB34A9375677541D749655CAAB779A26F826B57CE7203A22C24730D7099ADF";
   constant CPIX_NORMAL_INIT_53_BIT_13_C : bit_vector(255 downto 0) := x"42A2CE7EF1331DD5B7DCE511E323363670D7DC7FE72C73A6C0D3F98AC03D7628";
   constant CPIX_NORMAL_INIT_53_BIT_14_C : bit_vector(255 downto 0) := x"58D51CD12946FA82D7A72FE8A0789CD78B228EE2E2AF2D78C1148D3409706844";
   constant CPIX_NORMAL_INIT_54_BIT_00_C : bit_vector(255 downto 0) := x"5DA1EB7910EF1BC62809A60FD6C2616BD2139D58C4A581552CB518F5F5F14E96";
   constant CPIX_NORMAL_INIT_54_BIT_01_C : bit_vector(255 downto 0) := x"0ADF8C1BBC46EAD972C2517A4AEA9948FEE8C076E163CFE93C39B4F6409BFD13";
   constant CPIX_NORMAL_INIT_54_BIT_02_C : bit_vector(255 downto 0) := x"0B4D11988EC19D01C83E78E3D3D316A06E59B9079427F24BA581A7D9BE4EC200";
   constant CPIX_NORMAL_INIT_54_BIT_03_C : bit_vector(255 downto 0) := x"E273F690F3B6686846D20920AA45F44D76BDBF699332F4626CDA1F2BE34E8589";
   constant CPIX_NORMAL_INIT_54_BIT_04_C : bit_vector(255 downto 0) := x"533B800C3352D483FD2D683CF0406E586C7B4EFCB7130D9D903C3D6D753B1E1F";
   constant CPIX_NORMAL_INIT_54_BIT_05_C : bit_vector(255 downto 0) := x"7EB1466669393FC834C7ED1F4E1884B1AA29858DA49657FC2ED884B850799F1F";
   constant CPIX_NORMAL_INIT_54_BIT_06_C : bit_vector(255 downto 0) := x"F44E3FFAF70F41C54AAEEB1124DC19E7876D8F5B4DEB7DCD47B2CBE6218B5AFD";
   constant CPIX_NORMAL_INIT_54_BIT_07_C : bit_vector(255 downto 0) := x"B376536F4AA93A64012D32A35780DCC555C7ECF4C169873D365B1A0E8D938093";
   constant CPIX_NORMAL_INIT_54_BIT_08_C : bit_vector(255 downto 0) := x"DF57D99C3AA92D92EC552EB6A6AD2BBF69A0906167393A6FFCBE40C7ED75255B";
   constant CPIX_NORMAL_INIT_54_BIT_09_C : bit_vector(255 downto 0) := x"40A4BE259973EB3F80E74CC8EE177D896190CD676A9D254C31B3985466BBBDE9";
   constant CPIX_NORMAL_INIT_54_BIT_10_C : bit_vector(255 downto 0) := x"536155A1FF8F2535647C5C6981AF4F58D70F2AC61F83C27ED40A2BD044A70B19";
   constant CPIX_NORMAL_INIT_54_BIT_11_C : bit_vector(255 downto 0) := x"1258C1347C45BAEB24C06C90E05FA623419F3FC05CE6EC3E87C07EAD0108E793";
   constant CPIX_NORMAL_INIT_54_BIT_12_C : bit_vector(255 downto 0) := x"99EEEB1E239206DBCF8B3A486A251F7590B17BCDA78BCD30CB57DFD80E8C4433";
   constant CPIX_NORMAL_INIT_54_BIT_13_C : bit_vector(255 downto 0) := x"02FFE75ABB4C3C3811FCB0A2B31751AB3D4CFE05FC5114D4DC12B23392CA2AC3";
   constant CPIX_NORMAL_INIT_54_BIT_14_C : bit_vector(255 downto 0) := x"BB48D42B4016666026A40DE4D4CE1FF0F5482EBD06CDF6A869F5F6A7F462ED2F";
   constant CPIX_NORMAL_INIT_55_BIT_00_C : bit_vector(255 downto 0) := x"6740E8701183539E2E3720D048B905DE42DE32362A06EDBED79C1185BE173BF2";
   constant CPIX_NORMAL_INIT_55_BIT_01_C : bit_vector(255 downto 0) := x"35513B8D600C8FD15627860C365A1AD602F86F55D854D03BCC7C71F37DAA45C0";
   constant CPIX_NORMAL_INIT_55_BIT_02_C : bit_vector(255 downto 0) := x"0C252B6F16875C3F754E7106E31C33FA1763A33B0F0149039261580B40331240";
   constant CPIX_NORMAL_INIT_55_BIT_03_C : bit_vector(255 downto 0) := x"E10E407E5CE42A204E25673DDE00093940E034960200CAC6BA80741AFDCA2D05";
   constant CPIX_NORMAL_INIT_55_BIT_04_C : bit_vector(255 downto 0) := x"F2DB7AB7805B82450A1D8AFF4227B4DABB51130AFCBBD0B570E9828072F5ADFB";
   constant CPIX_NORMAL_INIT_55_BIT_05_C : bit_vector(255 downto 0) := x"D6F6807BC4BC6CABDA253FC603F6F173A3619C6F59F5EDC3B07C9723552E22BF";
   constant CPIX_NORMAL_INIT_55_BIT_06_C : bit_vector(255 downto 0) := x"D7533DF91330CD63E1721C7CAB974613FFA56A73D3FF75F38ED5072D175D645B";
   constant CPIX_NORMAL_INIT_55_BIT_07_C : bit_vector(255 downto 0) := x"C17377D7380B4A7DBF467D634551426F7F93CD71F7F72DBBED1859C9D257B873";
   constant CPIX_NORMAL_INIT_55_BIT_08_C : bit_vector(255 downto 0) := x"EE5059B210D37B1384844F6B4F7E3D362EBF056E34B7AB77FE9632174979A177";
   constant CPIX_NORMAL_INIT_55_BIT_09_C : bit_vector(255 downto 0) := x"64742591663D3927D39B504ED57D033C273DF8F67ABD7B6B09F7103D6534FA3D";
   constant CPIX_NORMAL_INIT_55_BIT_10_C : bit_vector(255 downto 0) := x"6E51534735DE531A38A344502F132C643DEE9270CA39F6A3DDD72956D0D28617";
   constant CPIX_NORMAL_INIT_55_BIT_11_C : bit_vector(255 downto 0) := x"41FDC69BD8CE89BC26ED172CD573771473861CFECA3D3385A69902317C824947";
   constant CPIX_NORMAL_INIT_55_BIT_12_C : bit_vector(255 downto 0) := x"4C9DA0EC3308076AB6CAA5D94BB4A0BC30C48762843D1BE9C663581FBD567E03";
   constant CPIX_NORMAL_INIT_55_BIT_13_C : bit_vector(255 downto 0) := x"6FCF47EA064F72860E78E3B271832500541826D4A235836536CAE8FDC9BAAB81";
   constant CPIX_NORMAL_INIT_55_BIT_14_C : bit_vector(255 downto 0) := x"24EC6A98335470A478CD79B776BF38D602E89FBA0E31406DC920048EC3187985";
   constant CPIX_NORMAL_INIT_56_BIT_00_C : bit_vector(255 downto 0) := x"E8B6BD3468F74F93C09AA28E91E38060252C5AE87C5538A3C00843A5B5C51736";
   constant CPIX_NORMAL_INIT_56_BIT_01_C : bit_vector(255 downto 0) := x"F05EBA655DCD3CC46797B4255B1F20517FA6B2E77ABA6D6BFDD8696508727263";
   constant CPIX_NORMAL_INIT_56_BIT_02_C : bit_vector(255 downto 0) := x"C6B88E71EF70D2297359A1D78484545EDF2DE9E12B084B3E04BED6496030BB24";
   constant CPIX_NORMAL_INIT_56_BIT_03_C : bit_vector(255 downto 0) := x"68251A122EB006B16F582FD1AA7D3C0D393D1FEC084D1A64E22BB8D7DD9A1A77";
   constant CPIX_NORMAL_INIT_56_BIT_04_C : bit_vector(255 downto 0) := x"E5AC1F36A8A338835C849890B9151297CD02C24AE27E433FD6938BC475A09030";
   constant CPIX_NORMAL_INIT_56_BIT_05_C : bit_vector(255 downto 0) := x"BDC3F4F00C52A84DCE13FF319980EAD604060CA9391147F4BF59E4C329FE669B";
   constant CPIX_NORMAL_INIT_56_BIT_06_C : bit_vector(255 downto 0) := x"397E86EB2999C17E46E95D8A4B33188C3EF8524BD2A969D9EF8C43902204E8D3";
   constant CPIX_NORMAL_INIT_56_BIT_07_C : bit_vector(255 downto 0) := x"BE1959BD4D86ABB6EB7FB5A36FBE8F3729A4E1D70D4F424BA744807A4719F557";
   constant CPIX_NORMAL_INIT_56_BIT_08_C : bit_vector(255 downto 0) := x"BE2AC94AD20A8F4407ACFF7741BADCFDCD4C9D1F4955153AA61D9741A2BD0D98";
   constant CPIX_NORMAL_INIT_56_BIT_09_C : bit_vector(255 downto 0) := x"DB8D8413BE25DA7F89C36C482DE41B30796B25EDE15DDDA10E828A1340D7FD22";
   constant CPIX_NORMAL_INIT_56_BIT_10_C : bit_vector(255 downto 0) := x"22F3F800327C26998D08C70C85C32688E8B8F75BAA2F08D5EC78DB0469D8E30C";
   constant CPIX_NORMAL_INIT_56_BIT_11_C : bit_vector(255 downto 0) := x"4E78E71CD992BF6DC8058955A47AF90C17E1CB65C75D28B321B923F9C821E56A";
   constant CPIX_NORMAL_INIT_56_BIT_12_C : bit_vector(255 downto 0) := x"1EF14DFA792C12BCFC944BC11587706F6B689A3570F1AF469E1400EC1AB9FD04";
   constant CPIX_NORMAL_INIT_56_BIT_13_C : bit_vector(255 downto 0) := x"EC445FF22D7FFE0A1FFAE0B39E9D2ABE695BA00FFCCA6CFD42B68723C60AA66C";
   constant CPIX_NORMAL_INIT_56_BIT_14_C : bit_vector(255 downto 0) := x"69B5980CB186598F6F7F3A8358F52B9325D7CF3EF213977344B3FE0E7BE921DA";
   constant CPIX_NORMAL_INIT_57_BIT_00_C : bit_vector(255 downto 0) := x"2F544311C90E40A473523226E7FBA6E200418E6710E4CA176969603330C133FE";
   constant CPIX_NORMAL_INIT_57_BIT_01_C : bit_vector(255 downto 0) := x"5166F276181AD79899204182011BCCF05A053FB97DD1A6972DD3A22AE6763712";
   constant CPIX_NORMAL_INIT_57_BIT_02_C : bit_vector(255 downto 0) := x"08137427015F6DEA0A29062473FC6C980113CB9A7CEC921BD7CDA47D31F2313C";
   constant CPIX_NORMAL_INIT_57_BIT_03_C : bit_vector(255 downto 0) := x"DD3E8345CAECD3712D547611A1574857AB4533E279B0EAA6A078077CE83D4445";
   constant CPIX_NORMAL_INIT_57_BIT_04_C : bit_vector(255 downto 0) := x"99DD0098B50FF8F9873DDA5E92D756D3D8EC888AEBE75977F44A7AFA8B24E92F";
   constant CPIX_NORMAL_INIT_57_BIT_05_C : bit_vector(255 downto 0) := x"D58163367D9D29BC7A80A46C47FFB3D5FFA6C942F03B1786099E51AEB0D4DADD";
   constant CPIX_NORMAL_INIT_57_BIT_06_C : bit_vector(255 downto 0) := x"53C303B9A5432E516237736D3977D64DA64F409D0E33C8CAF5A8F34B27106ED5";
   constant CPIX_NORMAL_INIT_57_BIT_07_C : bit_vector(255 downto 0) := x"3984A62F2BFD0EF1AF3743DB9321EF51C6759A4A02C21435C7047E9647BDFBA3";
   constant CPIX_NORMAL_INIT_57_BIT_08_C : bit_vector(255 downto 0) := x"37F27D94ED2722068145722D5EF70E70C8254A28170788D385FD56D3C44328BB";
   constant CPIX_NORMAL_INIT_57_BIT_09_C : bit_vector(255 downto 0) := x"6D50A1A2CD75E1ECE6DC43E1728B6809CD9C67DEE87F1B296A39D48922D241D7";
   constant CPIX_NORMAL_INIT_57_BIT_10_C : bit_vector(255 downto 0) := x"4534519E4D6BCE41A34B20F523AC497186F3810F3D87BF7A6DC364F9AC8D707E";
   constant CPIX_NORMAL_INIT_57_BIT_11_C : bit_vector(255 downto 0) := x"47EA28C73B59B123552401B0506F94197DC552CE7D8AF7BC96C49229D0BF734C";
   constant CPIX_NORMAL_INIT_57_BIT_12_C : bit_vector(255 downto 0) := x"692033627E4FFFC3167648CE79185F2ACCD3ACB76CE8722A8880477D0F7014F0";
   constant CPIX_NORMAL_INIT_57_BIT_13_C : bit_vector(255 downto 0) := x"23741D31F3641131050A271515F0DA7EC006CFF26F0C1BFB899F685A96024D12";
   constant CPIX_NORMAL_INIT_57_BIT_14_C : bit_vector(255 downto 0) := x"2A1225A83B165B668B92FE92924DF2A0C611483F29232D6E8973860AD47823C2";
   constant CPIX_NORMAL_INIT_58_BIT_00_C : bit_vector(255 downto 0) := x"5B04C4E0268AF2C2EB040C33765CE94D14F9E7E3FFC0096BA6EF4375C6558998";
   constant CPIX_NORMAL_INIT_58_BIT_01_C : bit_vector(255 downto 0) := x"220CCE7048F66B77FCC1A9F4346F141A77B7EB71D4661FCB7E0A9D07F20133C2";
   constant CPIX_NORMAL_INIT_58_BIT_02_C : bit_vector(255 downto 0) := x"9F97DE6D859C05FE563791D5EA945D2E4F1218ECED60A4B6FD0470E3C16AEF11";
   constant CPIX_NORMAL_INIT_58_BIT_03_C : bit_vector(255 downto 0) := x"5716E1DCF29528DDF7971AEC7CABE1929D69DD4B1CDE5E14E0367CC08585879D";
   constant CPIX_NORMAL_INIT_58_BIT_04_C : bit_vector(255 downto 0) := x"F3C985B0FA0D76BDF4849E3BF8C66D0507DBC341765FACC0DA44867666E3A884";
   constant CPIX_NORMAL_INIT_58_BIT_05_C : bit_vector(255 downto 0) := x"B6F51D7369455E033FF6C120DA646615CE1EFE2F3B9BD5D24979E7B87C17D455";
   constant CPIX_NORMAL_INIT_58_BIT_06_C : bit_vector(255 downto 0) := x"51BC71155A8C1B0A07288673FD2186AE4CB4C29648CCE1CAD19E18CA1DAD8ADB";
   constant CPIX_NORMAL_INIT_58_BIT_07_C : bit_vector(255 downto 0) := x"5210CBDB2186E7C81A080C82E3B3BC928FCCC13186A3B4CF351927432F89CFF5";
   constant CPIX_NORMAL_INIT_58_BIT_08_C : bit_vector(255 downto 0) := x"50DCC93C0A2B978B7889CDBD8DA420217A72C6D45493DF67AEE49F49D4E3BCC4";
   constant CPIX_NORMAL_INIT_58_BIT_09_C : bit_vector(255 downto 0) := x"2AA477D43C0E447A3E2078BA422F205FA3C48C8EDD8DC7FFD3535F670412CC36";
   constant CPIX_NORMAL_INIT_58_BIT_10_C : bit_vector(255 downto 0) := x"DD507F8AE1BFFE0CDBCF3451A6E22FCA4750B80FB9C75808533A62D580EA99EA";
   constant CPIX_NORMAL_INIT_58_BIT_11_C : bit_vector(255 downto 0) := x"6E3604613453BA8B8010AA97B399F4097B8610E2A614E6CB953E0F852796F612";
   constant CPIX_NORMAL_INIT_58_BIT_12_C : bit_vector(255 downto 0) := x"722791168E016D002828440ADB10B1AEAE673CB27ABDB20B3B5D99E9A0A0636C";
   constant CPIX_NORMAL_INIT_58_BIT_13_C : bit_vector(255 downto 0) := x"4B2CCC9090BBA7F41C008139E83006B151C24F1602AEFE7CDC920F92C99AF320";
   constant CPIX_NORMAL_INIT_58_BIT_14_C : bit_vector(255 downto 0) := x"07EA618ED65702DDF7D7F3F42EE8DDD8A79B9857B550DC6F4C70C84779CDDA1A";
   constant CPIX_NORMAL_INIT_59_BIT_00_C : bit_vector(255 downto 0) := x"2C3EAB836C1EDBA469275652957C72CA2FB91F204961CD09C25D720C7C940095";
   constant CPIX_NORMAL_INIT_59_BIT_01_C : bit_vector(255 downto 0) := x"542E6068C14B7C432F62FF07E6EBD6CAB2C40129056CC1217A0F02B692054586";
   constant CPIX_NORMAL_INIT_59_BIT_02_C : bit_vector(255 downto 0) := x"3A76C0C0D02436DD6165D4934468A57C05C566293E1F84F4A83205906F6B47AB";
   constant CPIX_NORMAL_INIT_59_BIT_03_C : bit_vector(255 downto 0) := x"A75C6F3666A5DA8376519F1D6080B18F22726A1A236847E5650544F5E722159C";
   constant CPIX_NORMAL_INIT_59_BIT_04_C : bit_vector(255 downto 0) := x"B9AD2D8C2C7A6DF4F7ACC252BEBED096939296966337EB7E4360DE97C027FF95";
   constant CPIX_NORMAL_INIT_59_BIT_05_C : bit_vector(255 downto 0) := x"0A401BABE026E9184A261FEAD114F609E2BF164F008F102181C66199B5290164";
   constant CPIX_NORMAL_INIT_59_BIT_06_C : bit_vector(255 downto 0) := x"4477951AB531B82E85C7A2BC0FCEBA15798B2614D0F2B0E1E15030C95B7714AF";
   constant CPIX_NORMAL_INIT_59_BIT_07_C : bit_vector(255 downto 0) := x"2E16B26F169663A075B6E26F9B41453DE288596FE526353163244AB20D20F0B7";
   constant CPIX_NORMAL_INIT_59_BIT_08_C : bit_vector(255 downto 0) := x"F3C2D18BEB0E9D24F8AFBDA5A6639B5149CC32AB4F49C5EB0269AB67A6B11AF6";
   constant CPIX_NORMAL_INIT_59_BIT_09_C : bit_vector(255 downto 0) := x"C71714476B5052BB209A2D2DB7B233ABD57AA20B0307BB05D9451FC7581622CD";
   constant CPIX_NORMAL_INIT_59_BIT_10_C : bit_vector(255 downto 0) := x"BD14D6801671B8405B1F83B7C9671CD5D636BC5CAC7C937324261AA695672765";
   constant CPIX_NORMAL_INIT_59_BIT_11_C : bit_vector(255 downto 0) := x"E043C7B7F31420297748F8FF23B0E96B1780E5176947D303E098DE2E969DCC93";
   constant CPIX_NORMAL_INIT_59_BIT_12_C : bit_vector(255 downto 0) := x"0F163CD96D36962C7C255A9446D1C3070DFB66A8D39FCCAD981273B7E3A8E9F8";
   constant CPIX_NORMAL_INIT_59_BIT_13_C : bit_vector(255 downto 0) := x"43F8188F6DABD2DF5A1284EAA604D9FF3F5D992E1B4ADCBE0DFA538A7311D92D";
   constant CPIX_NORMAL_INIT_59_BIT_14_C : bit_vector(255 downto 0) := x"06584521FD49C3335FCE79D944397772FB1D2876220F6CFD9C6927990F7B8C5F";
   constant CPIX_NORMAL_INIT_5A_BIT_00_C : bit_vector(255 downto 0) := x"5B00CCECB88BDEDC783E0270D8C23FFC7441C64B5B72C4BD54EA6A68E3766444";
   constant CPIX_NORMAL_INIT_5A_BIT_01_C : bit_vector(255 downto 0) := x"D2EB906C27B8DC24A52E5C9BF1E1561658522B2E175446603B69D57F9A765B34";
   constant CPIX_NORMAL_INIT_5A_BIT_02_C : bit_vector(255 downto 0) := x"8E43AF68152A559EC065A76D71BDE8D0BF833BDB74837079A7F7676EE02C7379";
   constant CPIX_NORMAL_INIT_5A_BIT_03_C : bit_vector(255 downto 0) := x"E0663F482F82764B928C1DFD9D69C5AC34FEF0D4A135BA8748FBB3EC81ABD563";
   constant CPIX_NORMAL_INIT_5A_BIT_04_C : bit_vector(255 downto 0) := x"84FD113130012BE876B9B040DC232C87B895B8894A636249A885023252C5EB5F";
   constant CPIX_NORMAL_INIT_5A_BIT_05_C : bit_vector(255 downto 0) := x"B0CED75244E3429FD1BD9177A2798603DE0DDE0970A4E1A49BD2DC32FDC983D8";
   constant CPIX_NORMAL_INIT_5A_BIT_06_C : bit_vector(255 downto 0) := x"66A6CD3A719CB8A1C94FBDE97CC0B4F66B28F2FF8C1F8831E0891C04748299E2";
   constant CPIX_NORMAL_INIT_5A_BIT_07_C : bit_vector(255 downto 0) := x"3AFABCBB87DF179976D3CD4DFA3842F529FC97DD5491951EBCCCD9BFC4B12791";
   constant CPIX_NORMAL_INIT_5A_BIT_08_C : bit_vector(255 downto 0) := x"C72E2D35DEB411A8973DD7B1C93B0B5143242CE31637D6BCF1ED55CEB9979145";
   constant CPIX_NORMAL_INIT_5A_BIT_09_C : bit_vector(255 downto 0) := x"10AC368D9B4240F509D29B42274C184C003CFBED9F3A6FEA0A6DF47DC2B58A8A";
   constant CPIX_NORMAL_INIT_5A_BIT_10_C : bit_vector(255 downto 0) := x"16C8D741CA263C22B74C6B578C06FF66B46E27E7FF626AB3E6DC0FF4542CF06C";
   constant CPIX_NORMAL_INIT_5A_BIT_11_C : bit_vector(255 downto 0) := x"D90436A6A604A92134A6DAA5830765A3FA944D4C07139A5855FFF2A7C0CA7560";
   constant CPIX_NORMAL_INIT_5A_BIT_12_C : bit_vector(255 downto 0) := x"3FD353289225A3880BC832D77FEA2CE9CE2FA5EBB6E607F365D3AA84AB94B9D1";
   constant CPIX_NORMAL_INIT_5A_BIT_13_C : bit_vector(255 downto 0) := x"88637B5D37DB54FEFFB42AC6F81D207FF48F5B529421B30B66961C163C357F5E";
   constant CPIX_NORMAL_INIT_5A_BIT_14_C : bit_vector(255 downto 0) := x"CFFA957305F37F79281DB81896862A3507E1FC001D7F23636A9478F7F04560D1";
   constant CPIX_NORMAL_INIT_5B_BIT_00_C : bit_vector(255 downto 0) := x"573098261073C978D475770D0EFDC3C66BD47CC87999C393898C5F5F7067C617";
   constant CPIX_NORMAL_INIT_5B_BIT_01_C : bit_vector(255 downto 0) := x"6A60DDD5F230868D214027AB702D3CBA1E1A48B44E3546F2338C2059289DDE33";
   constant CPIX_NORMAL_INIT_5B_BIT_02_C : bit_vector(255 downto 0) := x"4495CF9073126F76E037012066AF4BC2509146DA9A9D3301799C531099361F21";
   constant CPIX_NORMAL_INIT_5B_BIT_03_C : bit_vector(255 downto 0) := x"9ADED2C268B379CFBC4502AC2B91E039A5B8445D751D4064822DA91CD0D30863";
   constant CPIX_NORMAL_INIT_5B_BIT_04_C : bit_vector(255 downto 0) := x"F83A8B2B125C7FC8AACD0389C03BC7347A36AF6412980E3B04B1FEA69A26E49D";
   constant CPIX_NORMAL_INIT_5B_BIT_05_C : bit_vector(255 downto 0) := x"13573B29D3C228D9993195927197EAACEC0649086703A0D2B4F2F44083C8FD25";
   constant CPIX_NORMAL_INIT_5B_BIT_06_C : bit_vector(255 downto 0) := x"0ED3B845E3579990DA08079EF3F4DA7DCCBA404DD041B405516E640D0BB33152";
   constant CPIX_NORMAL_INIT_5B_BIT_07_C : bit_vector(255 downto 0) := x"52573DB08EA7588B2F6170ED5CB77541CD840D89DECA2112FE7894B1B69D8D3A";
   constant CPIX_NORMAL_INIT_5B_BIT_08_C : bit_vector(255 downto 0) := x"B27139922C98FA3635A03EED8D68DA1A9323F65AC8A69E14DC4E39BB0F00E7A4";
   constant CPIX_NORMAL_INIT_5B_BIT_09_C : bit_vector(255 downto 0) := x"5B2150B7928CDF85126289C6862128FF9AD9B3F22C782F8BDB4F7E36A59D93F5";
   constant CPIX_NORMAL_INIT_5B_BIT_10_C : bit_vector(255 downto 0) := x"667044B0779B84F99151D20688C262628C37663CADB77FA028F4C37636CF94E5";
   constant CPIX_NORMAL_INIT_5B_BIT_11_C : bit_vector(255 downto 0) := x"2962B716A55F74C23D56E359A281776E756B722B386D8E7478999739C738DB6F";
   constant CPIX_NORMAL_INIT_5B_BIT_12_C : bit_vector(255 downto 0) := x"2841DDDC1757208BC76491CB719716160D977AC3EABCDF68C62B6C78D819DB82";
   constant CPIX_NORMAL_INIT_5B_BIT_13_C : bit_vector(255 downto 0) := x"13FC33E0E32CCD2C0D21355B7B91087CA818338F6DB173D397D99D7886027E76";
   constant CPIX_NORMAL_INIT_5B_BIT_14_C : bit_vector(255 downto 0) := x"49B49ECB7637C9613CCFDEA24CEEB98E3C752EC9D60E879083C39C2DDEE8D113";
   constant CPIX_NORMAL_INIT_5C_BIT_00_C : bit_vector(255 downto 0) := x"2FFAB26BC59874C3AD7068CC2C3D2275A8112EA217828081445546F7739D753E";
   constant CPIX_NORMAL_INIT_5C_BIT_01_C : bit_vector(255 downto 0) := x"3FA900B8E434156EE185DB61B70F6B4360859465D4E4DC29B74CD0E43530BFA7";
   constant CPIX_NORMAL_INIT_5C_BIT_02_C : bit_vector(255 downto 0) := x"51D1FCF2E669DD1C0C862596ED49AFD15BA1EBBFF4AAA58424C00BBE6AB2115C";
   constant CPIX_NORMAL_INIT_5C_BIT_03_C : bit_vector(255 downto 0) := x"B01EA1E9123FD0E338D0E373030705C057605A008B607F1BAFDF8FEF47A9E703";
   constant CPIX_NORMAL_INIT_5C_BIT_04_C : bit_vector(255 downto 0) := x"DF97C740680CD2FC8BF9F292FFCD0294363CB83948CBC762BD38128BAC76B91D";
   constant CPIX_NORMAL_INIT_5C_BIT_05_C : bit_vector(255 downto 0) := x"A08EFAA7F92D5D1243C564A774C28FB032D98AA057396FEC97E932D4B7CB9DE1";
   constant CPIX_NORMAL_INIT_5C_BIT_06_C : bit_vector(255 downto 0) := x"9B5F47233890B68AFBFB2697ED7A00D76ADC69578A2D2E2CE1B67B527767452B";
   constant CPIX_NORMAL_INIT_5C_BIT_07_C : bit_vector(255 downto 0) := x"FD6685D78A0A2560CB155B163C4B9BF26DAC87331C5739C7D1579C355C3C289F";
   constant CPIX_NORMAL_INIT_5C_BIT_08_C : bit_vector(255 downto 0) := x"5AA429E1179FBD27E1CFCB505B858451DB60E18A0F806AD1CC34D006BE1D5AB9";
   constant CPIX_NORMAL_INIT_5C_BIT_09_C : bit_vector(255 downto 0) := x"679CF478E4B7FE2D99E92F0858CCB0E38C7EEA10FF21C47047CAE6EF7F832333";
   constant CPIX_NORMAL_INIT_5C_BIT_10_C : bit_vector(255 downto 0) := x"8B70D50DBB40A0B1477669801D7176A9B4BEFF6C5CE0FF0D4DFFCAE4C57D1BF8";
   constant CPIX_NORMAL_INIT_5C_BIT_11_C : bit_vector(255 downto 0) := x"FA05AF14354C03805E452CFC2CB4786BD52B06A69497537781FBAA712B2ADBE8";
   constant CPIX_NORMAL_INIT_5C_BIT_12_C : bit_vector(255 downto 0) := x"D02E9E2AD82024624728655F051FF38700C8F57F853FEE88682945CE5D9BEE0C";
   constant CPIX_NORMAL_INIT_5C_BIT_13_C : bit_vector(255 downto 0) := x"B84276EFF2417FD7EF58F0268D253C7AF02D0DF0AA2C20382DA6B767468BACF4";
   constant CPIX_NORMAL_INIT_5C_BIT_14_C : bit_vector(255 downto 0) := x"748E3CC123F7A4555EEE4B10A6E2BED4BF01E76ECB9178620A90689D3366CE98";
   constant CPIX_NORMAL_INIT_5D_BIT_00_C : bit_vector(255 downto 0) := x"644026CC4FE4E603166C795CA39C239922090CC813986D401B06FE5AA0E14795";
   constant CPIX_NORMAL_INIT_5D_BIT_01_C : bit_vector(255 downto 0) := x"50D4AD2D5F75D218178EEC4CE36883183244A238669AD79A4123108B2B1054EE";
   constant CPIX_NORMAL_INIT_5D_BIT_02_C : bit_vector(255 downto 0) := x"A165DC13E8C7CD9AFD9789A8EC9C8EBDC4826643A4BB3769AE79C584D6467786";
   constant CPIX_NORMAL_INIT_5D_BIT_03_C : bit_vector(255 downto 0) := x"1C3E5053432A2D84687BD62669FDD85C648C6DA961BD26A64778D4687613CDCD";
   constant CPIX_NORMAL_INIT_5D_BIT_04_C : bit_vector(255 downto 0) := x"F5C9704C9390376D96221871828C3CBCB84DE4718DD0EBFFDBA152F5839985C7";
   constant CPIX_NORMAL_INIT_5D_BIT_05_C : bit_vector(255 downto 0) := x"1D511F9B52F0A5BA51409AE3556A08F0362D744A70DB14FF0A21C5577820CF44";
   constant CPIX_NORMAL_INIT_5D_BIT_06_C : bit_vector(255 downto 0) := x"F0DEA1F2AFCC9FB10DCC6CC8568DB12F45DC99F844B7EAD3532830EA3B22F200";
   constant CPIX_NORMAL_INIT_5D_BIT_07_C : bit_vector(255 downto 0) := x"3F0CAF78EF3F2783146BF6DC45C8589A6442CA36318C683C628B2F2862FF89BB";
   constant CPIX_NORMAL_INIT_5D_BIT_08_C : bit_vector(255 downto 0) := x"79C872C68CD62D43274C9A1C68F0FC040449EBDB064263395A829AC8330FE077";
   constant CPIX_NORMAL_INIT_5D_BIT_09_C : bit_vector(255 downto 0) := x"3DACB98FDC85DB8C21BAC3FD1DC137701BFC94E02FB5153342E73C39085276C9";
   constant CPIX_NORMAL_INIT_5D_BIT_10_C : bit_vector(255 downto 0) := x"7AC0251A555540DB3042888B0860795B6A573DEB30A02F9938B1F59D2513563C";
   constant CPIX_NORMAL_INIT_5D_BIT_11_C : bit_vector(255 downto 0) := x"2175D7AF5F66258B25EF005A1D0E1318A377D32DFC6892961D3769DB3E39F9A6";
   constant CPIX_NORMAL_INIT_5D_BIT_12_C : bit_vector(255 downto 0) := x"170635841907CEFF543E5BC050F30D3D27347186FD34DC66C393CC5C86B8DEFE";
   constant CPIX_NORMAL_INIT_5D_BIT_13_C : bit_vector(255 downto 0) := x"794040084AA249B2B5CC7391F5FDA432093C3BF3E88EF98248671CB3D7DDDEF3";
   constant CPIX_NORMAL_INIT_5D_BIT_14_C : bit_vector(255 downto 0) := x"358487DE420788454B669C20AEBFD39342565847CAD6C2F106305FC9ADF89F1C";
   constant CPIX_NORMAL_INIT_5E_BIT_00_C : bit_vector(255 downto 0) := x"C3536691E32B2E36AE9188BCA21A4D30BD3C679B553736D176B8CD3CB572C656";
   constant CPIX_NORMAL_INIT_5E_BIT_01_C : bit_vector(255 downto 0) := x"0D7861121F0B3D13D2D95BFAEFF79D4D33957BB6D1F869642CFDE8D98EA457D9";
   constant CPIX_NORMAL_INIT_5E_BIT_02_C : bit_vector(255 downto 0) := x"9EC5EC5164AC34832546E7F598B8A15A8F5D2AFC35D80115DA7C4CAC4F705A02";
   constant CPIX_NORMAL_INIT_5E_BIT_03_C : bit_vector(255 downto 0) := x"4C58A18387916B60ABBDE37CA0016C07F8F0228ACDE69391026047263FA067D7";
   constant CPIX_NORMAL_INIT_5E_BIT_04_C : bit_vector(255 downto 0) := x"1806B77364D9F3C579E75430C78753B478E1E61FD52603D96269D9FCD32AA43D";
   constant CPIX_NORMAL_INIT_5E_BIT_05_C : bit_vector(255 downto 0) := x"679754BE70C48206761A256E813CD3CCA92EA755DD70B9DBD3F908F77B88E9AF";
   constant CPIX_NORMAL_INIT_5E_BIT_06_C : bit_vector(255 downto 0) := x"0F3AEE7060F9271FADB784F7CD5653EBAA1D1C8B05D8E51FF70745F20DCD7561";
   constant CPIX_NORMAL_INIT_5E_BIT_07_C : bit_vector(255 downto 0) := x"F2D87195EA5B43F543E8861959AB52DBD04768BB08F92C49931CB575E3652263";
   constant CPIX_NORMAL_INIT_5E_BIT_08_C : bit_vector(255 downto 0) := x"5CA48A8DA36EAD69871180F24E7C912563EBF71E59F52BB1EC84DB1A697FAE40";
   constant CPIX_NORMAL_INIT_5E_BIT_09_C : bit_vector(255 downto 0) := x"975CE912FDCD53ACEB0C88311B7644C9633FE8F2904212F72BF85808CCCEFC4B";
   constant CPIX_NORMAL_INIT_5E_BIT_10_C : bit_vector(255 downto 0) := x"F8766E73C50EB293A254048AF395CFAF6650685516F27588034EB2C723FD8023";
   constant CPIX_NORMAL_INIT_5E_BIT_11_C : bit_vector(255 downto 0) := x"870DC76940B2A16EAC06CC6B5ABF666EC18B4AE2A5BE9DD1128B09684C2D1EE9";
   constant CPIX_NORMAL_INIT_5E_BIT_12_C : bit_vector(255 downto 0) := x"E801E916E97FAF1A69E2B44A9966F77A65B9BE254C6198648F2559396A30DE92";
   constant CPIX_NORMAL_INIT_5E_BIT_13_C : bit_vector(255 downto 0) := x"2EC66FC98C60F6D20CB4EB354687ED41AA4741219F33448239AD9EF04BF7FD54";
   constant CPIX_NORMAL_INIT_5E_BIT_14_C : bit_vector(255 downto 0) := x"78CE9693BC0326F0B171FB3EF84F421E528F20F8E340B5ABBDDB2EB81C784C22";
   constant CPIX_NORMAL_INIT_5F_BIT_00_C : bit_vector(255 downto 0) := x"4E143B7D0B6D216443C648DDA2A7EAE75182FAAD64225FB623A644021690A946";
   constant CPIX_NORMAL_INIT_5F_BIT_01_C : bit_vector(255 downto 0) := x"12F63D981065D2C90604F725B666D6071B1C679F1F50A3CD0C7058C823D24971";
   constant CPIX_NORMAL_INIT_5F_BIT_02_C : bit_vector(255 downto 0) := x"EDA1922BE7B1438BD66A2B9C292F2463E02D9C03C9A40B29D87FFE30E17F2276";
   constant CPIX_NORMAL_INIT_5F_BIT_03_C : bit_vector(255 downto 0) := x"FFEB7DE7E61BF7C8779B00798F96C2DD1964B85A7FD3EB7E58ABC9F2559D3689";
   constant CPIX_NORMAL_INIT_5F_BIT_04_C : bit_vector(255 downto 0) := x"D22F562F53CDD53DA864E228962573ECB01FE969CE288797B2D9966DFB91762B";
   constant CPIX_NORMAL_INIT_5F_BIT_05_C : bit_vector(255 downto 0) := x"51E1E1071C6466EB217E60BD60534F7A2F91DFCB1265C7AF09B0BAC156D1F18E";
   constant CPIX_NORMAL_INIT_5F_BIT_06_C : bit_vector(255 downto 0) := x"418DC47957EA4A79228208711C355E2312F867EF6B80549D04DE9DDC652BA4E7";
   constant CPIX_NORMAL_INIT_5F_BIT_07_C : bit_vector(255 downto 0) := x"40B3D0E3DCE86F8C507A8598649E77DB201412175F17DD23A228D79AFDB10041";
   constant CPIX_NORMAL_INIT_5F_BIT_08_C : bit_vector(255 downto 0) := x"0A310B5F5DFD02D841BF530534210DEE3D5CF3EB2E30C193029C883284608B14";
   constant CPIX_NORMAL_INIT_5F_BIT_09_C : bit_vector(255 downto 0) := x"091651E30B0DCE6E50D80A2B3490E4FEF18E91238919A9A5777CC2AFB112D7A2";
   constant CPIX_NORMAL_INIT_5F_BIT_10_C : bit_vector(255 downto 0) := x"2DC66F89047F0FEC61AF66C3704995B06D0A95A9A132B05133A47736A5E00C25";
   constant CPIX_NORMAL_INIT_5F_BIT_11_C : bit_vector(255 downto 0) := x"0D84E39113BC507200F67A441144AB796A313A7FED8FDACF345548EB04364E99";
   constant CPIX_NORMAL_INIT_5F_BIT_12_C : bit_vector(255 downto 0) := x"05B036C16AF428CC245704DD411CA01E4FB739F6834211371BF3B13F1F2A2055";
   constant CPIX_NORMAL_INIT_5F_BIT_13_C : bit_vector(255 downto 0) := x"0490E01B099D230E0E6B77E76E1708291D7182FB49300FA20E67268504B5E461";
   constant CPIX_NORMAL_INIT_5F_BIT_14_C : bit_vector(255 downto 0) := x"003654104AA94CBAAE70C78BB0D69C8862FDF0974203C71447437C7967702F12";
   constant CPIX_NORMAL_INIT_60_BIT_00_C : bit_vector(255 downto 0) := x"5A3CCDD857B2753585A24E99A93DC3A1BF648DDC8FC1EF49DE26584DD0E990A6";
   constant CPIX_NORMAL_INIT_60_BIT_01_C : bit_vector(255 downto 0) := x"BEA4660B1F51E10B6596CCFE9DDD5E88286CDF6F517359FE11CE5380689737A9";
   constant CPIX_NORMAL_INIT_60_BIT_02_C : bit_vector(255 downto 0) := x"F40844B76A6ABDF6F1D0514D1B560B0ACEBB0E9DAF7EF279DBCFB30CB1A5A6DF";
   constant CPIX_NORMAL_INIT_60_BIT_03_C : bit_vector(255 downto 0) := x"18E533C4043FA9DE293C158ED3C4089F436A8BEF5C8283A95C50A9CEBA871FAF";
   constant CPIX_NORMAL_INIT_60_BIT_04_C : bit_vector(255 downto 0) := x"BE9B1A3CCB2AAF40D22341DA2D3B633433F06BF61BDC003D5CFC90DF96AAC1CE";
   constant CPIX_NORMAL_INIT_60_BIT_05_C : bit_vector(255 downto 0) := x"8A68BAAFC1BFB6233FDACF55FED5F60A075DF5E66E6BE5F1572FABACC109054B";
   constant CPIX_NORMAL_INIT_60_BIT_06_C : bit_vector(255 downto 0) := x"B04326EFD08F33FEE4E716CC35661E5A68E71D6914FAD9C17464F6D4FB419EDF";
   constant CPIX_NORMAL_INIT_60_BIT_07_C : bit_vector(255 downto 0) := x"69D725470EEB9C85E85427572B0A0C310030D71DD648F8031FE0FD775B9FC7AB";
   constant CPIX_NORMAL_INIT_60_BIT_08_C : bit_vector(255 downto 0) := x"52989F323B1E8344906DB13F67CEF8A759A7854A931482D11A359B065FC02D42";
   constant CPIX_NORMAL_INIT_60_BIT_09_C : bit_vector(255 downto 0) := x"F96F6A9F638B861F2B09DDB9E1F08377C824874CC0A5AE5659081BC62C39477E";
   constant CPIX_NORMAL_INIT_60_BIT_10_C : bit_vector(255 downto 0) := x"C36BE435E4B7185229B286D6538705431884C466931872961EA3D2071F9C3CBC";
   constant CPIX_NORMAL_INIT_60_BIT_11_C : bit_vector(255 downto 0) := x"BC058BE16E319F3A6C0C7F199ACC23A5267AEDBF12C90F52131BAF106A61A49C";
   constant CPIX_NORMAL_INIT_60_BIT_12_C : bit_vector(255 downto 0) := x"847FB87FC367D9AFB64DF04B1718F6C736FE46247A52CEEC05D08855239A75C4";
   constant CPIX_NORMAL_INIT_60_BIT_13_C : bit_vector(255 downto 0) := x"318FF108340FA6D84EC8D1FDF6A1063A57E0324D160334383FB70E7B0C368CC0";
   constant CPIX_NORMAL_INIT_60_BIT_14_C : bit_vector(255 downto 0) := x"49E0332ACD71EA46DDCA1248A1A60BB12FF3B021336E5F25B3A5D8F22EE95070";
   constant CPIX_NORMAL_INIT_61_BIT_00_C : bit_vector(255 downto 0) := x"EE6D4B625739B6EF9F94CB7D97F0E6FD7B557B5B9388C8AE6C64D8A5675C1011";
   constant CPIX_NORMAL_INIT_61_BIT_01_C : bit_vector(255 downto 0) := x"508C5CC00382D0A466CB6FCC50EAB31080BA5A353EC9F4471796026C0A97E560";
   constant CPIX_NORMAL_INIT_61_BIT_02_C : bit_vector(255 downto 0) := x"867B38A6309C83EFBFB56033B6033DA362FF14236262299290FF901D2F7DD94B";
   constant CPIX_NORMAL_INIT_61_BIT_03_C : bit_vector(255 downto 0) := x"5B61903C8719FA7B3B018D6306B61E937709FC8C3E33BDFE41673436FEA18DF6";
   constant CPIX_NORMAL_INIT_61_BIT_04_C : bit_vector(255 downto 0) := x"22EC803A5F65B8DF192E7A3B660068E585B54C566CA591B1501CDE60F72E4C02";
   constant CPIX_NORMAL_INIT_61_BIT_05_C : bit_vector(255 downto 0) := x"77001AFB0CED5FDA3F5BDB302BF031F7E83D7713912DF03575AF6CC33943AAB0";
   constant CPIX_NORMAL_INIT_61_BIT_06_C : bit_vector(255 downto 0) := x"EBE6F6A47813014673A8AA1E34EBEB30A94A7E0A7704F1C6BFFE492F71A03E7C";
   constant CPIX_NORMAL_INIT_61_BIT_07_C : bit_vector(255 downto 0) := x"5A4E345F19E8F9623D0684E3685B82039A64017A5AFA4675B471AB2A99069D3F";
   constant CPIX_NORMAL_INIT_61_BIT_08_C : bit_vector(255 downto 0) := x"4BB315F8031BE854718887361147AD0063A7258EFCC9C0599D4D9D9D6D3E0F99";
   constant CPIX_NORMAL_INIT_61_BIT_09_C : bit_vector(255 downto 0) := x"58BEE8995546AFA6364A7D683664D3DC9B4B930D7466BFA5DF0ECF99971BD3D7";
   constant CPIX_NORMAL_INIT_61_BIT_10_C : bit_vector(255 downto 0) := x"61660D55036F8C2256D77A6642CE5F7BDA1FFC899FCCA3FD238F764CE0C2DC4C";
   constant CPIX_NORMAL_INIT_61_BIT_11_C : bit_vector(255 downto 0) := x"07B51C3D584409B646EFC24ADBF0EE76DEB067F02A8DA7E475DA4FDA5984B01B";
   constant CPIX_NORMAL_INIT_61_BIT_12_C : bit_vector(255 downto 0) := x"7096BF3C475C6171A459FBC0D23940560977B8745C1B190B3A77E474C222FA31";
   constant CPIX_NORMAL_INIT_61_BIT_13_C : bit_vector(255 downto 0) := x"410102A9DF62649607E8F7D588AF675CCECC0A1A3CDAF7BEB9335B1CE5FF7F2A";
   constant CPIX_NORMAL_INIT_61_BIT_14_C : bit_vector(255 downto 0) := x"50F48531BEE5D23D328DF8CEA1C14571F43743CD63C90CC87B4DF1A2275255B3";
   constant CPIX_NORMAL_INIT_62_BIT_00_C : bit_vector(255 downto 0) := x"9F7E1E5D86E0E9E040AA77AE0ED3483FC1F363F2AF2F97AEF99E96ABE7625B85";
   constant CPIX_NORMAL_INIT_62_BIT_01_C : bit_vector(255 downto 0) := x"48C8C65B267F9594C769E95222801037DF081A19B4654A6A355E90F795B6AF4B";
   constant CPIX_NORMAL_INIT_62_BIT_02_C : bit_vector(255 downto 0) := x"D4183A74F93DC77AE8B7B42442DEECAD3507177E7F35307B05C0F201CADB814A";
   constant CPIX_NORMAL_INIT_62_BIT_03_C : bit_vector(255 downto 0) := x"50D60C535EE76BF6928BBC95C879DE4C236BB706B2541717777DC58336A93266";
   constant CPIX_NORMAL_INIT_62_BIT_04_C : bit_vector(255 downto 0) := x"323A80643EE0016D1E8F7F5C93755B1B1F0F548879A00BFA059E3705E420E771";
   constant CPIX_NORMAL_INIT_62_BIT_05_C : bit_vector(255 downto 0) := x"E556F47BDDB383921148AA27EE90A462B13F1238A734074E2732CB50666F8969";
   constant CPIX_NORMAL_INIT_62_BIT_06_C : bit_vector(255 downto 0) := x"4A45E8F9CA10B604D8A087988BB7A0DB5D5DD7E946904E0D90C0E7BCB21A5910";
   constant CPIX_NORMAL_INIT_62_BIT_07_C : bit_vector(255 downto 0) := x"60ED39D6AEEA10084C26B58E34A2869EB930463F12F3201F52331D0C5087EE7A";
   constant CPIX_NORMAL_INIT_62_BIT_08_C : bit_vector(255 downto 0) := x"495DFC689A029E8BB30CD1A1543DB16918A29F05B6F8A708CE9EE422A81CCCA7";
   constant CPIX_NORMAL_INIT_62_BIT_09_C : bit_vector(255 downto 0) := x"22D71B7A26724A0AE53D9260DCF59896CB22E43440927515081E6EE621E15575";
   constant CPIX_NORMAL_INIT_62_BIT_10_C : bit_vector(255 downto 0) := x"D1AFF8B7B3AE55BD6AD3CBA0C509CC45F25AE75AD71662326CF4553D770AF05E";
   constant CPIX_NORMAL_INIT_62_BIT_11_C : bit_vector(255 downto 0) := x"3200EC62EC03A440DA9CF0F6B0A343BF7077E43FFCE9FAC379FB8FC6E002B623";
   constant CPIX_NORMAL_INIT_62_BIT_12_C : bit_vector(255 downto 0) := x"66741008E0B6180A6D8C2B826E22523A1F839EF5AACF666856D9A4C112105D7C";
   constant CPIX_NORMAL_INIT_62_BIT_13_C : bit_vector(255 downto 0) := x"2AC9B3E082C08E08D0ECE2ED2A5B30A57D3CDA2C641D68EC60A0CF121EF14CC5";
   constant CPIX_NORMAL_INIT_62_BIT_14_C : bit_vector(255 downto 0) := x"3BB72D713BCDE3F71339E89FD139C5E6EC7A1F323F783C0879CF7341DD651640";
   constant CPIX_NORMAL_INIT_63_BIT_00_C : bit_vector(255 downto 0) := x"8DC7749FC04A83AE77824BCCB31AA620AADE61925CECD45EB5BF8456332664F2";
   constant CPIX_NORMAL_INIT_63_BIT_01_C : bit_vector(255 downto 0) := x"51E53723715F4257E03F42E97A045BB7141FAD39404EF4AFD0A90B2EF6C050AC";
   constant CPIX_NORMAL_INIT_63_BIT_02_C : bit_vector(255 downto 0) := x"36D5BB27300D3E734005C26EE8E73989B5CE5DE7295630F68D56F15652EC3029";
   constant CPIX_NORMAL_INIT_63_BIT_03_C : bit_vector(255 downto 0) := x"E9A94DAB2AE32A1AA61E33F158111D861BF3E6560C24E0E9EADC9A8D3832F233";
   constant CPIX_NORMAL_INIT_63_BIT_04_C : bit_vector(255 downto 0) := x"35D386EF75AAD365E10467C793974CC47B75D2D61881D66581FDEBD6BB70B02F";
   constant CPIX_NORMAL_INIT_63_BIT_05_C : bit_vector(255 downto 0) := x"50DD8B0A353103293207B543A77544BFC77C5045C54406894F895F94AC81419D";
   constant CPIX_NORMAL_INIT_63_BIT_06_C : bit_vector(255 downto 0) := x"25CB427DD2793B286B1760AF4607496D2987D63C50AC54828C07981FE08A9ABE";
   constant CPIX_NORMAL_INIT_63_BIT_07_C : bit_vector(255 downto 0) := x"650F4EB046274C2EDBC4BAD1FB635C990AD088C596C6CA9A751C2F5F1DC4DEE6";
   constant CPIX_NORMAL_INIT_63_BIT_08_C : bit_vector(255 downto 0) := x"E7EFE0CA9B497FA6D9EA920D8059B92422AAFA74C4145997FEC52D79F2841631";
   constant CPIX_NORMAL_INIT_63_BIT_09_C : bit_vector(255 downto 0) := x"66F0F490B6FA8100ED7BE7D71BAFE3C80A9F3B68A6A8DF18012C4106E1D17C90";
   constant CPIX_NORMAL_INIT_63_BIT_10_C : bit_vector(255 downto 0) := x"33C19FE78123E0440375D7B3968E3A78DBB6262F5A1333D3F97FF338A22AF580";
   constant CPIX_NORMAL_INIT_63_BIT_11_C : bit_vector(255 downto 0) := x"03765176A437AD7E4C44EF444F586E27E01DE9648907E6F552991634B00E721D";
   constant CPIX_NORMAL_INIT_63_BIT_12_C : bit_vector(255 downto 0) := x"05DD0C744470CD15BE4BE049AA0D65FCBEA637B2A0CEA0E729F21FAFE6866AEE";
   constant CPIX_NORMAL_INIT_63_BIT_13_C : bit_vector(255 downto 0) := x"6B869A1764585D0CFD4C732016E76C4ADC6DEC00567F50F3F2BA0F5B7DF16D28";
   constant CPIX_NORMAL_INIT_63_BIT_14_C : bit_vector(255 downto 0) := x"02A887731BBEF2BAA518C489F8C43D5A370B277CC5C347DB0C4A26B0174FD7ED";
   constant CPIX_NORMAL_INIT_64_BIT_00_C : bit_vector(255 downto 0) := x"D76620D6458977AF67F708B88C0CD7E06B5FB9AAB62381EE868400001E45ABE9";
   constant CPIX_NORMAL_INIT_64_BIT_01_C : bit_vector(255 downto 0) := x"582623E9D95BC8A0135FD90547461C6F0750338F711B7A10DE3374986311D863";
   constant CPIX_NORMAL_INIT_64_BIT_02_C : bit_vector(255 downto 0) := x"F5CBA4DE6C9D77A9E04EEF3FAC3ACF10BFDB51E9455EB9D4466C06F4C45A1BA5";
   constant CPIX_NORMAL_INIT_64_BIT_03_C : bit_vector(255 downto 0) := x"23EC53A502C2E7DDE1A465646BDE4B65B5DC27452AB20655CF6540AA2CE5DD56";
   constant CPIX_NORMAL_INIT_64_BIT_04_C : bit_vector(255 downto 0) := x"23720A37E3F206807323B570E66E659191AC64F80C14AFD3375F1C564827E1E1";
   constant CPIX_NORMAL_INIT_64_BIT_05_C : bit_vector(255 downto 0) := x"BC4E06A3F50E69DE833EA881E0C4BE2732BD01096EB6FA030E088722BD3C8184";
   constant CPIX_NORMAL_INIT_64_BIT_06_C : bit_vector(255 downto 0) := x"131A4AC9C7AB44C60C93264E8FC19EC1E5617491EDB10DB5824FCD4F38DABB77";
   constant CPIX_NORMAL_INIT_64_BIT_07_C : bit_vector(255 downto 0) := x"01B0C6F30A7A89404DAE943CCA71829E2AE075EB26B4CA6A377BC2E6B4F52F51";
   constant CPIX_NORMAL_INIT_64_BIT_08_C : bit_vector(255 downto 0) := x"C8262C364FFC7243BA78D4F1D1DE09FB1ED84570587B6C69CC03D0B215F5CD36";
   constant CPIX_NORMAL_INIT_64_BIT_09_C : bit_vector(255 downto 0) := x"7123BCE7E380690DAE87FD91BFAE6175EFA9B6CE2CED65FC467606F8510C1B87";
   constant CPIX_NORMAL_INIT_64_BIT_10_C : bit_vector(255 downto 0) := x"28B4696E029AE93EA8677A9EF0D425BADC4FEF2385B627F10E9C27F18B90A50F";
   constant CPIX_NORMAL_INIT_64_BIT_11_C : bit_vector(255 downto 0) := x"119CA2A456A350CCDBED1FDA24D6995C948F0FBEFA415969F9229BE0368122BB";
   constant CPIX_NORMAL_INIT_64_BIT_12_C : bit_vector(255 downto 0) := x"786D74200003E87AADFDA4D712B7CBD73BD20ABBFCF832A2535078A971575EA2";
   constant CPIX_NORMAL_INIT_64_BIT_13_C : bit_vector(255 downto 0) := x"26A0D9EDD37338528581EE599CE6B452457962178E03C8E1F9477227C6DCBBA1";
   constant CPIX_NORMAL_INIT_64_BIT_14_C : bit_vector(255 downto 0) := x"126D1B60693E7EA90ED6ABDD50E5BA8DA2A81BB3031B9255F68ED54201AB55D9";
   constant CPIX_NORMAL_INIT_65_BIT_00_C : bit_vector(255 downto 0) := x"803659FFF855BA6D8E4551D9A6D266EA834050A3891A866BD9E473AB886836AF";
   constant CPIX_NORMAL_INIT_65_BIT_01_C : bit_vector(255 downto 0) := x"4F68B30B6C31B27B55B13D349F214BBC117B3C989E4B609D04FBF976B541D754";
   constant CPIX_NORMAL_INIT_65_BIT_02_C : bit_vector(255 downto 0) := x"56BB0359A40080C72DBE0B53E8080646AAD31C73475FCE51ADE2634BB7ADCF8B";
   constant CPIX_NORMAL_INIT_65_BIT_03_C : bit_vector(255 downto 0) := x"AC98A27E30DF8158255E7CD204178CB126D621316918878C7F4A63FF9DEAE3A7";
   constant CPIX_NORMAL_INIT_65_BIT_04_C : bit_vector(255 downto 0) := x"56AD6439B96142DA344383527A4559B60BDAC8BB40399FF75B74BC9BA9E97714";
   constant CPIX_NORMAL_INIT_65_BIT_05_C : bit_vector(255 downto 0) := x"355ACC78F2D5177B20AF61940542D9D7A442ECECF44E597DA265EAC0CC428E67";
   constant CPIX_NORMAL_INIT_65_BIT_06_C : bit_vector(255 downto 0) := x"6757DE671EA05653A496C736EA410F8231E94CA89597E2F8F2B980465582AAA3";
   constant CPIX_NORMAL_INIT_65_BIT_07_C : bit_vector(255 downto 0) := x"33360414FE84D2A64BED7C6BA93215BF59DEA70B4EF803DAAC59498384C382E9";
   constant CPIX_NORMAL_INIT_65_BIT_08_C : bit_vector(255 downto 0) := x"23A29A4939A0312A2E5BEC741632167FE36E9DDD8FE89E2B31A2252F7D64785D";
   constant CPIX_NORMAL_INIT_65_BIT_09_C : bit_vector(255 downto 0) := x"1309A103A375F4BE12364234C6847877A8846659E2824753F43190B5CED88D61";
   constant CPIX_NORMAL_INIT_65_BIT_10_C : bit_vector(255 downto 0) := x"F5C765B060574BFAF0F3DBEEE1EBD780B0BE1F48A7997DAA12C100B5815908B5";
   constant CPIX_NORMAL_INIT_65_BIT_11_C : bit_vector(255 downto 0) := x"802BCD337A2A6EE07996696948C7E13F89B8D2A14F4A2D7D3FCFEE5B4A8A0C31";
   constant CPIX_NORMAL_INIT_65_BIT_12_C : bit_vector(255 downto 0) := x"CC8215E9D9B75E77699C83F8FAD034C039E7CA199C6B19377DE6D12636F6FF8F";
   constant CPIX_NORMAL_INIT_65_BIT_13_C : bit_vector(255 downto 0) := x"8E9FFB350B075B4F1C2F38AF2698595C4E63FA37E9C850F85D6117E034DBFB1C";
   constant CPIX_NORMAL_INIT_65_BIT_14_C : bit_vector(255 downto 0) := x"5D1F701FC60FDBC16EF6F2E0EB1FABB8449608DC82645FF74D549D62D515F565";
   constant CPIX_NORMAL_INIT_66_BIT_00_C : bit_vector(255 downto 0) := x"A9B09E4F0ED843F5E927CF3869AB269ED68D65C50B11BB2AC93DE636BB0A7CF8";
   constant CPIX_NORMAL_INIT_66_BIT_01_C : bit_vector(255 downto 0) := x"7B27CC8ADA2BF7A9482AE42611D95AEA022D5463AE6B038C40D278AB4C39EF41";
   constant CPIX_NORMAL_INIT_66_BIT_02_C : bit_vector(255 downto 0) := x"298CF5B8C4844F7B8216B0FB5027454A5E348E14568408516F376A1774BD2F1E";
   constant CPIX_NORMAL_INIT_66_BIT_03_C : bit_vector(255 downto 0) := x"A3830BF7841302E10DEC9C3764237FD222B0A108D91E1C8A26570F49534A0B37";
   constant CPIX_NORMAL_INIT_66_BIT_04_C : bit_vector(255 downto 0) := x"95AF2B991FB4F5E025E18398892344951B99391498111F7CC30726CE72EF991C";
   constant CPIX_NORMAL_INIT_66_BIT_05_C : bit_vector(255 downto 0) := x"E79E52D6267469521C217FD999F6D89EBDA1ACC9C2E3E92E25B9E13AE84416ED";
   constant CPIX_NORMAL_INIT_66_BIT_06_C : bit_vector(255 downto 0) := x"586007A71F88C5F9369C6C3E16BDFD80EEEA7FF5FD6237F4825914F402694F69";
   constant CPIX_NORMAL_INIT_66_BIT_07_C : bit_vector(255 downto 0) := x"E335610976992754793884F48F74D3357CCD36F7656A4C6BF12E2F454C19756D";
   constant CPIX_NORMAL_INIT_66_BIT_08_C : bit_vector(255 downto 0) := x"F5DD108AB8FE331BDAB11D4F3E1A878F36B487F20F7664DB902D527D456F4243";
   constant CPIX_NORMAL_INIT_66_BIT_09_C : bit_vector(255 downto 0) := x"021AAE6CB48F18B04658DFE32C1697C73E7B6FDB125B4EFCEC312A553E3E1453";
   constant CPIX_NORMAL_INIT_66_BIT_10_C : bit_vector(255 downto 0) := x"678516BF8E4D5F53D8CE2CB1747121355B40F649C17001FD4641136E5965654B";
   constant CPIX_NORMAL_INIT_66_BIT_11_C : bit_vector(255 downto 0) := x"6955EF1B8D221082B19BB404537B71F560F86459503D26C23F147065C9DCBCD5";
   constant CPIX_NORMAL_INIT_66_BIT_12_C : bit_vector(255 downto 0) := x"CB7F3DE6265C69ADA5CD1698BC4D6DC041246F50D12B4C21F9C68ADD68248BD9";
   constant CPIX_NORMAL_INIT_66_BIT_13_C : bit_vector(255 downto 0) := x"2F675A1EE4A5C2D4D06225A0D5D0F41E58D2A7528A8E8FA23BE710A73DB33BBF";
   constant CPIX_NORMAL_INIT_66_BIT_14_C : bit_vector(255 downto 0) := x"E9213371D9CC139207B39E233D833E072BEC0F48A89F180D4DFF41F361932892";
   constant CPIX_NORMAL_INIT_67_BIT_00_C : bit_vector(255 downto 0) := x"CEBAFDC2405D9D98F09C947DBC8648FFE576B9A42A8BD9FE774D7C5BF8122D04";
   constant CPIX_NORMAL_INIT_67_BIT_01_C : bit_vector(255 downto 0) := x"7236FA55B36B626B1A411BF1168BC919683B59B0D65721CEBCA086D95A773588";
   constant CPIX_NORMAL_INIT_67_BIT_02_C : bit_vector(255 downto 0) := x"05721B5C674B320CF8702AE41A109E64EC0F2C45033EFBF16DE458B4B68975B2";
   constant CPIX_NORMAL_INIT_67_BIT_03_C : bit_vector(255 downto 0) := x"DA15E7B98DF9745E8E56555903DB431E5C1C6112D878C12339DC5D5A33C0E25A";
   constant CPIX_NORMAL_INIT_67_BIT_04_C : bit_vector(255 downto 0) := x"323F30C91A1E16AB271471E118A257666D5ED384ADBF5A1EAF359BA179558D69";
   constant CPIX_NORMAL_INIT_67_BIT_05_C : bit_vector(255 downto 0) := x"E6483A1625C88D202EA19C33D636D6D97DD6E2CAA65CCF501B7A3A2D684F5EC6";
   constant CPIX_NORMAL_INIT_67_BIT_06_C : bit_vector(255 downto 0) := x"47CC052647196B53FC27256726AB5A721677CD0184F76A8F349D524C6430B33E";
   constant CPIX_NORMAL_INIT_67_BIT_07_C : bit_vector(255 downto 0) := x"423A37DEE6472D7E94FBE6F42152BB1106A1ED3CB863C116AFB6A4FF70FE4E4A";
   constant CPIX_NORMAL_INIT_67_BIT_08_C : bit_vector(255 downto 0) := x"71D7203F77486E149BE10E0174EA38199D7C9A5D2ECCB5523A6FDFE5881C892A";
   constant CPIX_NORMAL_INIT_67_BIT_09_C : bit_vector(255 downto 0) := x"11A68B5D6C0B27D32E8105E28F0E29DD4B965657052FA4A8850B629EF679949D";
   constant CPIX_NORMAL_INIT_67_BIT_10_C : bit_vector(255 downto 0) := x"12F5B52D2A4D072615C34B9A546C8CE08A67053A0917E04B981538A46BC2C0E2";
   constant CPIX_NORMAL_INIT_67_BIT_11_C : bit_vector(255 downto 0) := x"3BBAC64E4F400215F10069F158D7699F771D065586272FC6845CC862C01EB849";
   constant CPIX_NORMAL_INIT_67_BIT_12_C : bit_vector(255 downto 0) := x"0226F53B482D09708055534C1B2396E92B58B1C36E1F0B58D08D4FB44AD01BC8";
   constant CPIX_NORMAL_INIT_67_BIT_13_C : bit_vector(255 downto 0) := x"234C4617537934248C6B102038ECB3310D321FABB812B6F17BE32AD81F2B731B";
   constant CPIX_NORMAL_INIT_67_BIT_14_C : bit_vector(255 downto 0) := x"2086637EED83F0EC87202141063E0E41157DF7636FE6F8E13FAA24D9C0BDC8DF";
   constant CPIX_NORMAL_INIT_68_BIT_00_C : bit_vector(255 downto 0) := x"C9C3E96AB7969296695CFC5A8712BA287F1482B7CB196D7CC596CF2067E48BE0";
   constant CPIX_NORMAL_INIT_68_BIT_01_C : bit_vector(255 downto 0) := x"994A8F021843A5FC44F838FCB6626AAC6F126FE99686B8259E1CC1ACD5C63899";
   constant CPIX_NORMAL_INIT_68_BIT_02_C : bit_vector(255 downto 0) := x"9423BB0ED6A335FA969D825EEC8BAAE3859D9A540DCDDC50405616CEC340756F";
   constant CPIX_NORMAL_INIT_68_BIT_03_C : bit_vector(255 downto 0) := x"0BBA7ABFB4A31C901D1B691EFCE4E29ACEA4A02B1264771D7CCA019C6BC502BF";
   constant CPIX_NORMAL_INIT_68_BIT_04_C : bit_vector(255 downto 0) := x"B2D450AC1198296A22A4A0F723AD1DDA7FEB24D4D9F8054D98179498657997D3";
   constant CPIX_NORMAL_INIT_68_BIT_05_C : bit_vector(255 downto 0) := x"1C4F12BB1B616E1995C117C048ADC83C57DB79E9DB007665BF2AC4F8BDC5B0C4";
   constant CPIX_NORMAL_INIT_68_BIT_06_C : bit_vector(255 downto 0) := x"157062EE3600BE0F8405FF00E018478C4FBBEBCAD8AE4A1230ED902039BE88FC";
   constant CPIX_NORMAL_INIT_68_BIT_07_C : bit_vector(255 downto 0) := x"5C5393289980B70C33039AC31EFB7733BBC8C148FEB14CAB0A78CF967A0D0EAF";
   constant CPIX_NORMAL_INIT_68_BIT_08_C : bit_vector(255 downto 0) := x"1DDD26A73134530FA905654117E697DAB617520138496111FCE70EEAE5C68FAF";
   constant CPIX_NORMAL_INIT_68_BIT_09_C : bit_vector(255 downto 0) := x"4CA45098AB9095019133A58E0555172595EAAE3AD0938BA1FA8E1475D604B4DE";
   constant CPIX_NORMAL_INIT_68_BIT_10_C : bit_vector(255 downto 0) := x"B9580B583D6779C6C88CD17FF9D96FEE092BE9266C9A9F409179060EEB7AD5AC";
   constant CPIX_NORMAL_INIT_68_BIT_11_C : bit_vector(255 downto 0) := x"C1E547EBDF7F5FF5F1D1225E7A5CA553170246EE5F6C74F6C33D2FED215A2EE4";
   constant CPIX_NORMAL_INIT_68_BIT_12_C : bit_vector(255 downto 0) := x"EB58AD69D56FCA599E509E9E7AACADECFEB6145F52CF43C8125B32A7534BE2E1";
   constant CPIX_NORMAL_INIT_68_BIT_13_C : bit_vector(255 downto 0) := x"A7FA05DE746F6F52226B55AE4AE7E95AA297116A42978F4547D357B7AD61DB3A";
   constant CPIX_NORMAL_INIT_68_BIT_14_C : bit_vector(255 downto 0) := x"2BF072781EE7CD662FB7D6665F5909D593D1C0066382C3CB69DCAC0ADF6FC401";
   constant CPIX_NORMAL_INIT_69_BIT_00_C : bit_vector(255 downto 0) := x"AB9F2784C50A80411F666B926B88DC53E5C5D8116D35483E9FECCB241C5FBD23";
   constant CPIX_NORMAL_INIT_69_BIT_01_C : bit_vector(255 downto 0) := x"BA3C83F958BED5E7F3EF81EA7BA9EE899D3C54AA701C549F1C95F22D920FFF1D";
   constant CPIX_NORMAL_INIT_69_BIT_02_C : bit_vector(255 downto 0) := x"B7120B9F3D8F48E34487AC8A775BEFE925D4AE5B5B2107B38C5321DE026F1A8B";
   constant CPIX_NORMAL_INIT_69_BIT_03_C : bit_vector(255 downto 0) := x"609259809F1FBD8A99AB14977365D95638BD8927E8DD694D9B3F767493900919";
   constant CPIX_NORMAL_INIT_69_BIT_04_C : bit_vector(255 downto 0) := x"D6369CAEBA01297716C5D04C5068346BAB2CB89221D26AB5EBF64A1AA12AF02F";
   constant CPIX_NORMAL_INIT_69_BIT_05_C : bit_vector(255 downto 0) := x"1560B1F022449585DD959910C800344FE7318C20F07E25AA51FE4C6FF8B28F62";
   constant CPIX_NORMAL_INIT_69_BIT_06_C : bit_vector(255 downto 0) := x"4917307B8854348299BD2C189FD5F19D14267B6A40411DBD1EA6568C2E9DE6E5";
   constant CPIX_NORMAL_INIT_69_BIT_07_C : bit_vector(255 downto 0) := x"04FEFA8931D5998C768DEF11F7853F8F294D4FE09A8BCEA778CD2F054AA9B1B8";
   constant CPIX_NORMAL_INIT_69_BIT_08_C : bit_vector(255 downto 0) := x"41A2009BAEF40D80263C1528B5786275CAC1415EC63D2779FF0B4178BE711980";
   constant CPIX_NORMAL_INIT_69_BIT_09_C : bit_vector(255 downto 0) := x"486628A40CD1790CF73BFED5B95A532B10C1DBDB227BD41C0150377F975C18B2";
   constant CPIX_NORMAL_INIT_69_BIT_10_C : bit_vector(255 downto 0) := x"F0B9AF8E67BC9F3C82F447D7995CA9DF131B7773E5924C7AEB50381EDAD76C5F";
   constant CPIX_NORMAL_INIT_69_BIT_11_C : bit_vector(255 downto 0) := x"79551C9A92430DCEA168FB67A50AF78260AE8FF5AE690C5BB6EB98DAC7A97E4E";
   constant CPIX_NORMAL_INIT_69_BIT_12_C : bit_vector(255 downto 0) := x"5F4E51502490BF5B5E5C6D47591492BB7AB78558739A6150CCA6055BFB3BCCF1";
   constant CPIX_NORMAL_INIT_69_BIT_13_C : bit_vector(255 downto 0) := x"1DB7C528DAC0D55549A7D65D89EB8656540D2DA24232A4C152B1C2DFE88C32FF";
   constant CPIX_NORMAL_INIT_69_BIT_14_C : bit_vector(255 downto 0) := x"282861F99D7EC6A9B5BDDF6680A4246024A3112F2B5713F72ADE00996F5C2CDF";
   constant CPIX_NORMAL_INIT_6A_BIT_00_C : bit_vector(255 downto 0) := x"AF1BF6E48AB7D1F4E4AA8E1065F70E82D309F0C69D2C66B86E5D737F93D333C6";
   constant CPIX_NORMAL_INIT_6A_BIT_01_C : bit_vector(255 downto 0) := x"EF61B45C9F2582CDFADA2E97C3BA618AE8AA113CC42B591A90D8B6C1F51E3827";
   constant CPIX_NORMAL_INIT_6A_BIT_02_C : bit_vector(255 downto 0) := x"8B76AD63C964529BF55D3E31D5910592F202A8A42345D90472B9B79259C8C396";
   constant CPIX_NORMAL_INIT_6A_BIT_03_C : bit_vector(255 downto 0) := x"48078834BC72B0A6EC411EA9B9D3EBE215D8DD621924B0C25EEEA7C57A37D38C";
   constant CPIX_NORMAL_INIT_6A_BIT_04_C : bit_vector(255 downto 0) := x"D37D0390BA9F154B1013E18C4F085C6D17825189E666C0726736F32A96664737";
   constant CPIX_NORMAL_INIT_6A_BIT_05_C : bit_vector(255 downto 0) := x"9D878E6F3C791DC5D4A72CE9C795075F7C15667A49E3328CF68AEB1E6A8E06B7";
   constant CPIX_NORMAL_INIT_6A_BIT_06_C : bit_vector(255 downto 0) := x"916E14A5CD26F911FC759F4DB9161243C37FD3083FF04A2D96B30D6A1DBD4B3A";
   constant CPIX_NORMAL_INIT_6A_BIT_07_C : bit_vector(255 downto 0) := x"85596336F965001779A4DD6FE32A91E5D5173E74065D18A809EC86965333A989";
   constant CPIX_NORMAL_INIT_6A_BIT_08_C : bit_vector(255 downto 0) := x"F02D0971803737657F074DF5F85126C5B1AA7E69E07DDE7F6C845677EF09E443";
   constant CPIX_NORMAL_INIT_6A_BIT_09_C : bit_vector(255 downto 0) := x"444856659B03861656ED7E772D0644F60CF4A5F78D2AF16A48A57A424DA05FEE";
   constant CPIX_NORMAL_INIT_6A_BIT_10_C : bit_vector(255 downto 0) := x"70114B136D0071646F94B6DDA9618991140CFB4446268F329379399783780D32";
   constant CPIX_NORMAL_INIT_6A_BIT_11_C : bit_vector(255 downto 0) := x"0E9BABAE5E168550592FB658DA146921128460FF4868C3D50B782DE7987E02D9";
   constant CPIX_NORMAL_INIT_6A_BIT_12_C : bit_vector(255 downto 0) := x"2ACE5217DBCA3CCE4895863E9523E171AFF3591BBB7274348C7ADBA4B1BA3A05";
   constant CPIX_NORMAL_INIT_6A_BIT_13_C : bit_vector(255 downto 0) := x"7B1F135936DD49400258D4945BEEAFF81FD3F2660ECDD10F62F0E008A1D59B79";
   constant CPIX_NORMAL_INIT_6A_BIT_14_C : bit_vector(255 downto 0) := x"4E7A504C6A6D5F691EBF3406A40B9268F28701545C2C8B3CC27E1ADE6CDDC5E7";
   constant CPIX_NORMAL_INIT_6B_BIT_00_C : bit_vector(255 downto 0) := x"8FEF5CF3AEAA2022FF4AF34E99BAB7A0121B92C67424727BB9C19F927DE337EA";
   constant CPIX_NORMAL_INIT_6B_BIT_01_C : bit_vector(255 downto 0) := x"8A3A7F690AA3238ECF349B97F06D62F1D1EFB8AE2DE0413BC41CE0F5978712BF";
   constant CPIX_NORMAL_INIT_6B_BIT_02_C : bit_vector(255 downto 0) := x"AB6F5F0E3CB67E68CEBBFD950AEE6FE68EBF641076E9C83836ECF2A71A11565E";
   constant CPIX_NORMAL_INIT_6B_BIT_03_C : bit_vector(255 downto 0) := x"2DBAE29468F2E1213E5DFDF9C63EC4A0643A7C1C5658B65A663EA2B4C7E8B93F";
   constant CPIX_NORMAL_INIT_6B_BIT_04_C : bit_vector(255 downto 0) := x"A22083EE9E11B919A0AB6C25C357B447CE3FED692CA8E001A193579799B85C8E";
   constant CPIX_NORMAL_INIT_6B_BIT_05_C : bit_vector(255 downto 0) := x"88756A6E70C63FD8FDA1C7192B0FC8BAE9C621E2B5F4A8F9012E609CF2C97F51";
   constant CPIX_NORMAL_INIT_6B_BIT_06_C : bit_vector(255 downto 0) := x"193EC17055564592D30A35ABCED35078679D6A871A2B352A7E139EEAFA1840E9";
   constant CPIX_NORMAL_INIT_6B_BIT_07_C : bit_vector(255 downto 0) := x"68F77E3CF51B94F094B3190490791EFDF22E29FDF7CD7FB56CC92393D08712C1";
   constant CPIX_NORMAL_INIT_6B_BIT_08_C : bit_vector(255 downto 0) := x"5D48E55180563D34A43611A98E19816FF7A393B01EF50FAEA2A32087D290DE2A";
   constant CPIX_NORMAL_INIT_6B_BIT_09_C : bit_vector(255 downto 0) := x"60CDA4CEDA1C5B62AA5BE736768A5909BA81F4B7A9626C34674EC22C39B109E5";
   constant CPIX_NORMAL_INIT_6B_BIT_10_C : bit_vector(255 downto 0) := x"040B27B0D34C5E249D8369F7694EEA475DE0565AA292895AEED3F728E6B06AD2";
   constant CPIX_NORMAL_INIT_6B_BIT_11_C : bit_vector(255 downto 0) := x"1F6972C5040C0782681B6BDE98968F5236D2A9F6A0A0C7E21CB4926D4E5EA4C7";
   constant CPIX_NORMAL_INIT_6B_BIT_12_C : bit_vector(255 downto 0) := x"645573F9152B6237A9ED6E57A816340C3C2F661EE838094776B44CF1B00E3EE0";
   constant CPIX_NORMAL_INIT_6B_BIT_13_C : bit_vector(255 downto 0) := x"5424D40403500CB781BD723FAB639121E03D67F33FCDBA7F63C3EB6E1D9593D6";
   constant CPIX_NORMAL_INIT_6B_BIT_14_C : bit_vector(255 downto 0) := x"714E7135B9F992DC90276567A59386596CA2C92B77792C7949B7D1950DF37E4B";
   constant CPIX_NORMAL_INIT_6C_BIT_00_C : bit_vector(255 downto 0) := x"98069C439AEE79A481CBDB5D6DAD97F7CF73A4260FDAAD1DF12207D820EB6F55";
   constant CPIX_NORMAL_INIT_6C_BIT_01_C : bit_vector(255 downto 0) := x"9F401F22EF1FA63F59CDDDD91EB007FE9DC78953E736EA1EACD682E3534ABF0C";
   constant CPIX_NORMAL_INIT_6C_BIT_02_C : bit_vector(255 downto 0) := x"ED889858CE8726E2099FAAD5E9A870E934F50A0D129A503B912CE60DE007A8F4";
   constant CPIX_NORMAL_INIT_6C_BIT_03_C : bit_vector(255 downto 0) := x"5A7544B9DAB468EB54FADE4D48ACD5EA158BD86ADB2C6FD126A32930C56AA09E";
   constant CPIX_NORMAL_INIT_6C_BIT_04_C : bit_vector(255 downto 0) := x"E66A676C5495DFA99911DDB61C198518DE8DF25ECAB7E9701B9053E8B0977DEC";
   constant CPIX_NORMAL_INIT_6C_BIT_05_C : bit_vector(255 downto 0) := x"303FC5E2353B80F2DF138304814AC604D82460317F84B440B3F77B8926DC4184";
   constant CPIX_NORMAL_INIT_6C_BIT_06_C : bit_vector(255 downto 0) := x"0583C4E789DE3BD06B500DCCC04A350F0E403A331495E49F2C992ACB8B2B2EBF";
   constant CPIX_NORMAL_INIT_6C_BIT_07_C : bit_vector(255 downto 0) := x"71D7195C4DD7B006DA27C544543D24CD10BB49DA3229DDE9BA849DCB42517AB8";
   constant CPIX_NORMAL_INIT_6C_BIT_08_C : bit_vector(255 downto 0) := x"D98BF3A4EFECD5B02A5F328F16F5DC3D0AA6379B6AAEAC44759809B5FCB28DE8";
   constant CPIX_NORMAL_INIT_6C_BIT_09_C : bit_vector(255 downto 0) := x"9101701F4B66DD5F87D311F0A039215A7C586307746F1743D8ABAA9F913501A5";
   constant CPIX_NORMAL_INIT_6C_BIT_10_C : bit_vector(255 downto 0) := x"E09814E0339DA52895E2E695453D8554A07BCFF2BB40DD7B10E3E92217588FAF";
   constant CPIX_NORMAL_INIT_6C_BIT_11_C : bit_vector(255 downto 0) := x"C19DD04652EF5CE718C16191CAB79AA9750441FB80F9DAC2790DD0DB873859D1";
   constant CPIX_NORMAL_INIT_6C_BIT_12_C : bit_vector(255 downto 0) := x"316A6596643818912F5E9BAEA15DDEEE5581B0606603B0CFF56D7ED372AECC56";
   constant CPIX_NORMAL_INIT_6C_BIT_13_C : bit_vector(255 downto 0) := x"1E2B6F9B318FD0AF72A733AF2F1B50A636A88FDC2086E41C09311FF6A939ABD4";
   constant CPIX_NORMAL_INIT_6C_BIT_14_C : bit_vector(255 downto 0) := x"1204E2953B6A0655F265536EA65A37A31F4B911AD9DC7EAADBA1C0A724A16AB3";
   constant CPIX_NORMAL_INIT_6D_BIT_00_C : bit_vector(255 downto 0) := x"EB5AFA597BADC1668795956655CCBA6ECF51144598EB5681BF6CCA71F0892ABF";
   constant CPIX_NORMAL_INIT_6D_BIT_01_C : bit_vector(255 downto 0) := x"9FF22EC33BF28709B4B9A17B0F8ED0DB50D74AE15FC09A909E1BDA65860E9F8B";
   constant CPIX_NORMAL_INIT_6D_BIT_02_C : bit_vector(255 downto 0) := x"83EA7B34FEA4DE398C8A3B326F9C357EF1A7074A9C165C68677383275D5FCCDD";
   constant CPIX_NORMAL_INIT_6D_BIT_03_C : bit_vector(255 downto 0) := x"38DB476BDABEF8C64A824326936E996F85737913822EB68E49C846D82FD6870C";
   constant CPIX_NORMAL_INIT_6D_BIT_04_C : bit_vector(255 downto 0) := x"E7F5107AE0BA079475741B150DF1A5808E05407E5EC0B569E8EA3752E81518FB";
   constant CPIX_NORMAL_INIT_6D_BIT_05_C : bit_vector(255 downto 0) := x"1136996AA42949FEE12250C9CCC09AE4CB900D1B8E85C691B2B24ECCB9A5EA92";
   constant CPIX_NORMAL_INIT_6D_BIT_06_C : bit_vector(255 downto 0) := x"39E0D1A8B23BDCB6AF0280C007423D415DA74AECA3EE68CD76DFA1A4CA2049AD";
   constant CPIX_NORMAL_INIT_6D_BIT_07_C : bit_vector(255 downto 0) := x"116CBD2B746E2D40A82ABB41F68CDAA77FEF9B1A59A2F61C6E9A0883EAAF8C58";
   constant CPIX_NORMAL_INIT_6D_BIT_08_C : bit_vector(255 downto 0) := x"D4696AF54C5EA6B395D3ADB0A36F30DC9764BC0E969CA730146D159ECE0BE980";
   constant CPIX_NORMAL_INIT_6D_BIT_09_C : bit_vector(255 downto 0) := x"340D9AB815A9946FBADD667BB375CA9C0E5AB10C29B1522206FEB77F36C69CBB";
   constant CPIX_NORMAL_INIT_6D_BIT_10_C : bit_vector(255 downto 0) := x"540C5B8E8091A955A556ED7C6C955B8C1A90B565D271A1F5C75DF57DDA3C06C6";
   constant CPIX_NORMAL_INIT_6D_BIT_11_C : bit_vector(255 downto 0) := x"65D1C34961D2D857475766B46A9696B7A05DD0E44DBC914DF82211B20FDD8B44";
   constant CPIX_NORMAL_INIT_6D_BIT_12_C : bit_vector(255 downto 0) := x"60AA114B948B49112979FEB69766A2B9791694DA3A597F6EB7CFDD1D49F8F8E8";
   constant CPIX_NORMAL_INIT_6D_BIT_13_C : bit_vector(255 downto 0) := x"1E5CD6A624437826E25B6C599AA69175A5725B0FFC79E247CB3184D359216473";
   constant CPIX_NORMAL_INIT_6D_BIT_14_C : bit_vector(255 downto 0) := x"2CBB55A46BBD2FEB647A939899A6BE81BF850D7662E299741CE02755786DC048";
   constant CPIX_NORMAL_INIT_6E_BIT_00_C : bit_vector(255 downto 0) := x"BFA5C32EE99D25A5ADD5E59FCE0C33E7802875B61B9599AB1F82E677FFE2A5B8";
   constant CPIX_NORMAL_INIT_6E_BIT_01_C : bit_vector(255 downto 0) := x"B743F7BCF27FF337FD03BE04CB0743E8FE26B1B1D3214ADA57066AD12D6EE145";
   constant CPIX_NORMAL_INIT_6E_BIT_02_C : bit_vector(255 downto 0) := x"73A02A8709B3CB9B24506B523C8C92B988CDE7123A48EA722BFDAD99655DDC02";
   constant CPIX_NORMAL_INIT_6E_BIT_03_C : bit_vector(255 downto 0) := x"1401156C67846FA36E6E6E5D1E82530A43CE369D7AD5190A17309462DEFF9ED1";
   constant CPIX_NORMAL_INIT_6E_BIT_04_C : bit_vector(255 downto 0) := x"DA42985295249B6FC6C488FFB41C9889B990428EACD9F21A55E62B95E25B65E2";
   constant CPIX_NORMAL_INIT_6E_BIT_05_C : bit_vector(255 downto 0) := x"303B1CCF00BD062D52434B0F348164B0CBFDE621184D49BE5BBC167E9E18DBAC";
   constant CPIX_NORMAL_INIT_6E_BIT_06_C : bit_vector(255 downto 0) := x"DBCDFABC2A6A1AC60AAE0DF9164F75D0B31568DBFF59E70B7B61B676CD715507";
   constant CPIX_NORMAL_INIT_6E_BIT_07_C : bit_vector(255 downto 0) := x"62F6F75907DA0A2B41B54A665B765FAFE589B344B03163BF6F95216981A4266B";
   constant CPIX_NORMAL_INIT_6E_BIT_08_C : bit_vector(255 downto 0) := x"6A59A96152B26CE002FB115639BA53C53C6C1BE5CBB03882B5CB3878A481F23E";
   constant CPIX_NORMAL_INIT_6E_BIT_09_C : bit_vector(255 downto 0) := x"6EEBA8BA4F9E28543E8C7C051D66215A5AC6CDF6AE722ACFA6F0F4841BDF7955";
   constant CPIX_NORMAL_INIT_6E_BIT_10_C : bit_vector(255 downto 0) := x"7843000B41AB2463716F4C7A6CCA4116B482F0CC1568245CCFF62CF22FBC863E";
   constant CPIX_NORMAL_INIT_6E_BIT_11_C : bit_vector(255 downto 0) := x"449F354B4F032312D596E699256B76EDF0F04218306E6C67871D89158FF477BE";
   constant CPIX_NORMAL_INIT_6E_BIT_12_C : bit_vector(255 downto 0) := x"114821BF07380D265449E4A599A29EBF87B7A445164303D90AC787FA660B2BF2";
   constant CPIX_NORMAL_INIT_6E_BIT_13_C : bit_vector(255 downto 0) := x"60023D2DCA58CEC5267DEBE9252D9ABDE15FD079F2C5A467C62CF6466DD51BEC";
   constant CPIX_NORMAL_INIT_6E_BIT_14_C : bit_vector(255 downto 0) := x"489B11A035A4FF991121B99C143AEEB24B685DC03F30DDF8F0D7B865386A55BA";
   constant CPIX_NORMAL_INIT_6F_BIT_00_C : bit_vector(255 downto 0) := x"CF89C9BBE6D52202F601BAC2A2FEE71E6EA7288A07512CDB19A4FAA7A1593A6E";
   constant CPIX_NORMAL_INIT_6F_BIT_01_C : bit_vector(255 downto 0) := x"D2E3CD21F601F793C45A8A1886D4BE3A48E61BEB9D6ED17941D974C3CFB38674";
   constant CPIX_NORMAL_INIT_6F_BIT_02_C : bit_vector(255 downto 0) := x"2E16153A717B454702A126362520614FF04646C3449CAE9AB3FE3A83373F3655";
   constant CPIX_NORMAL_INIT_6F_BIT_03_C : bit_vector(255 downto 0) := x"FD6DD2FA3B07B99824E37BF72FAD2A5062CF98F6FAD6C079EDDB9D1B15047E1D";
   constant CPIX_NORMAL_INIT_6F_BIT_04_C : bit_vector(255 downto 0) := x"97171AA6C4D7945EC3E6B499DA96D85761D34A5A6D0499046D53951957AE95C2";
   constant CPIX_NORMAL_INIT_6F_BIT_05_C : bit_vector(255 downto 0) := x"0CC1247F474F413778BB149F2CF818CB190D48935347869AE6D0B4EA9F2D7AEF";
   constant CPIX_NORMAL_INIT_6F_BIT_06_C : bit_vector(255 downto 0) := x"0A861F16592524351E5F780A0BAA47CD37F44E51ED8DA11FF22B1AC3D00D2A44";
   constant CPIX_NORMAL_INIT_6F_BIT_07_C : bit_vector(255 downto 0) := x"0D8DAE7A078B4B5B401131A5D69BEC00DA48F31C1E922F1B816F3E6292C4D455";
   constant CPIX_NORMAL_INIT_6F_BIT_08_C : bit_vector(255 downto 0) := x"34332E1A0F11442F62DF74891AA584B02CBAD7E6908D36845FD33C7CE8B367F0";
   constant CPIX_NORMAL_INIT_6F_BIT_09_C : bit_vector(255 downto 0) := x"210D32B70A3648CFCB85A2EC569FC19D92E1EA1EF2A4350A57ED911D7E22ABE3";
   constant CPIX_NORMAL_INIT_6F_BIT_10_C : bit_vector(255 downto 0) := x"697A073E4F59428C638EC5C05C55CC24E57583D9D00BD8BF50600D4A13D95E85";
   constant CPIX_NORMAL_INIT_6F_BIT_11_C : bit_vector(255 downto 0) := x"28D81E050D7000F67477EBBB402F053A92960DC7E1A73F578B3DCFA81B26263E";
   constant CPIX_NORMAL_INIT_6F_BIT_12_C : bit_vector(255 downto 0) := x"0C587C6A410A02C33D6D91053DC73740E0E1E7F36DC3A5D74EF424A4B42674B9";
   constant CPIX_NORMAL_INIT_6F_BIT_13_C : bit_vector(255 downto 0) := x"08C32A53375D7126249F243D35580CC4797AA4D92CF419E0F104B5096EBC3DE0";
   constant CPIX_NORMAL_INIT_6F_BIT_14_C : bit_vector(255 downto 0) := x"05003E2FF49BC9AA5EC91190116654716B99E15CC4F7E3131B4ED0CFEB7E2625";
   constant CPIX_NORMAL_INIT_70_BIT_00_C : bit_vector(255 downto 0) := x"09CAE920474963218F8C65509B53ADFFC955E2BB72C519630B55470D4ADD7172";
   constant CPIX_NORMAL_INIT_70_BIT_01_C : bit_vector(255 downto 0) := x"03E2F0AC1C336CF100B81F918245943B3506D2783B6AB3596DE2422241C5182C";
   constant CPIX_NORMAL_INIT_70_BIT_02_C : bit_vector(255 downto 0) := x"96AFAABFF844B14C5F8D50790DC3F298C309B5D5FA422072B67AB5D6FB17DCFB";
   constant CPIX_NORMAL_INIT_70_BIT_03_C : bit_vector(255 downto 0) := x"340432D770A53D39526275FF05047CB52D5887FB544B986B17FF299E60EEE91F";
   constant CPIX_NORMAL_INIT_70_BIT_04_C : bit_vector(255 downto 0) := x"5E8714EB2777706C8C216C9C02B4D731FA3637E0854B67145C3D3A066E8F9F8B";
   constant CPIX_NORMAL_INIT_70_BIT_05_C : bit_vector(255 downto 0) := x"503F2E3B73B45C4DE65186D44F6961ECB6FF8FD57BF0F8D312CD77CC57FA8203";
   constant CPIX_NORMAL_INIT_70_BIT_06_C : bit_vector(255 downto 0) := x"FDDC61015EF34FF4E37350D9FF274C76C15F8B5FCD5A45336D260FA804D8F0BB";
   constant CPIX_NORMAL_INIT_70_BIT_07_C : bit_vector(255 downto 0) := x"33432EE5618D6391B4073F04C4F7A1A769413FA8E0117324049292E13CE53B9F";
   constant CPIX_NORMAL_INIT_70_BIT_08_C : bit_vector(255 downto 0) := x"3D0E13E04A9501E05D4BEA82A2AA673A1AB5739086C75BED2D83909834B13861";
   constant CPIX_NORMAL_INIT_70_BIT_09_C : bit_vector(255 downto 0) := x"2FEA01FD5366549AB39245FCB3BA9399E77B5B9372AECC95A4928CF122396617";
   constant CPIX_NORMAL_INIT_70_BIT_10_C : bit_vector(255 downto 0) := x"452017A519751B37B3EABADE5B52C9A297C4CD216D991901288592593D913A6E";
   constant CPIX_NORMAL_INIT_70_BIT_11_C : bit_vector(255 downto 0) := x"1C26202D1F93BCF5BC5C7ADC4B3B28C3E0BC74B76272BA5C57EF1A3113F074CA";
   constant CPIX_NORMAL_INIT_70_BIT_12_C : bit_vector(255 downto 0) := x"49F61244C2F8960125E4232375C495F487E795AFD2C312D95F1471BE08A05B48";
   constant CPIX_NORMAL_INIT_70_BIT_13_C : bit_vector(255 downto 0) := x"001EB5491ED8AF52BA336BDFE532CF774BC243DA3A8EDC171C5211467D3725A8";
   constant CPIX_NORMAL_INIT_70_BIT_14_C : bit_vector(255 downto 0) := x"0C84FC965AEBC804C51A5A2A72CD510D2C57A4F1AB12CD3C7DC45734DCAD7E04";
   constant CPIX_NORMAL_INIT_71_BIT_00_C : bit_vector(255 downto 0) := x"56B47C60A6C52C2B04B6D17C307EAAB248CD6313F0A0C6D872A2086014602AC7";
   constant CPIX_NORMAL_INIT_71_BIT_01_C : bit_vector(255 downto 0) := x"5AE13F7161DB5C160750D2B3BE4972BC625E349B66419EDDC090CC5757EDA734";
   constant CPIX_NORMAL_INIT_71_BIT_02_C : bit_vector(255 downto 0) := x"0A557E152056E168CF3DB17D91893CF6C238C6848DC49D3601977C071CB09987";
   constant CPIX_NORMAL_INIT_71_BIT_03_C : bit_vector(255 downto 0) := x"EC2F4173F31C202939C1B4FEEAB2456549293D7D9BE822A25751D81142A95E51";
   constant CPIX_NORMAL_INIT_71_BIT_04_C : bit_vector(255 downto 0) := x"499F4F94E05999287499B8A48EF9F4E7178C7C063B729433330A643F0B70C4D4";
   constant CPIX_NORMAL_INIT_71_BIT_05_C : bit_vector(255 downto 0) := x"0AB3441671C1D40F9600103A3A38E82AC1CFAD9902F5F8C5C716D413559057A6";
   constant CPIX_NORMAL_INIT_71_BIT_06_C : bit_vector(255 downto 0) := x"4B169676514F112669961E29A1A3CB9F30E6B0D0AC9ABDCB229E183288DED320";
   constant CPIX_NORMAL_INIT_71_BIT_07_C : bit_vector(255 downto 0) := x"433C1527B8F8F52A38A8899B427328BD4E69FF0225CB4D9BE4171D43152209F7";
   constant CPIX_NORMAL_INIT_71_BIT_08_C : bit_vector(255 downto 0) := x"DFCBB27DAF9282E45FF48029F866D81422E6B1BBD28C06C62DB0DED2BBC5E2AD";
   constant CPIX_NORMAL_INIT_71_BIT_09_C : bit_vector(255 downto 0) := x"5CC8DF80E7D93FDA3B76DEB20601C86859375533C694ACA9B5C40940237D4C04";
   constant CPIX_NORMAL_INIT_71_BIT_10_C : bit_vector(255 downto 0) := x"58BD85C0149D9B76BD573159E7D6D7C88FEDDF0E79BC82A0D3D391556C0653C3";
   constant CPIX_NORMAL_INIT_71_BIT_11_C : bit_vector(255 downto 0) := x"1505C5E720F03275C2E4A1DC1A14C35250E5E1C0BACDCD1F45C7EEF96FB9C1D5";
   constant CPIX_NORMAL_INIT_71_BIT_12_C : bit_vector(255 downto 0) := x"0A2404A0F3C2F24EFD5DCBCD6D3FD97F5402CD236A79751739BCFB561AC81026";
   constant CPIX_NORMAL_INIT_71_BIT_13_C : bit_vector(255 downto 0) := x"79B14222E2541D63A6E0170DDF336C667ADC98B28EDE734C66B6426E4CB13C28";
   constant CPIX_NORMAL_INIT_71_BIT_14_C : bit_vector(255 downto 0) := x"1E953FDFC28AE8635356891B235C139E7D647ADD16EB868DE73576626B50A410";
   constant CPIX_NORMAL_INIT_72_BIT_00_C : bit_vector(255 downto 0) := x"7AD01F094FF526A06FF25C6853A059A06AB6F5A0A2D15D638C102A7067FFCF01";
   constant CPIX_NORMAL_INIT_72_BIT_01_C : bit_vector(255 downto 0) := x"4C037BDE4391929E6898EF225C4599304FE8560CB1714C449C4B6900D2B59FA4";
   constant CPIX_NORMAL_INIT_72_BIT_02_C : bit_vector(255 downto 0) := x"5712DB812CA0E09191B55F90BD53C79B816B3E5E63A6ABF0770E2BE854A90C3C";
   constant CPIX_NORMAL_INIT_72_BIT_03_C : bit_vector(255 downto 0) := x"AAD7508243E9012C59D42E9A635FAEDD5E3C0DDAEC447374CE505510F4AE60A1";
   constant CPIX_NORMAL_INIT_72_BIT_04_C : bit_vector(255 downto 0) := x"1E46F41B4111702D3B3F0ABD34EBEE505515D91875C4D7088A4E20F9138125CC";
   constant CPIX_NORMAL_INIT_72_BIT_05_C : bit_vector(255 downto 0) := x"43A6C8174F4801A9C1FECB26D4F8A1B5E31DC36BB7E8C8F55E027DF13215E688";
   constant CPIX_NORMAL_INIT_72_BIT_06_C : bit_vector(255 downto 0) := x"51B53C11C995F0394E3E81DEDE8109FD133A9F090953B8B8C448EC2C93A36BF5";
   constant CPIX_NORMAL_INIT_72_BIT_07_C : bit_vector(255 downto 0) := x"5500F89D3E67E50F2BC33E1BE229899E0C9D37A02F86B49B7C4F5CB7579DCC70";
   constant CPIX_NORMAL_INIT_72_BIT_08_C : bit_vector(255 downto 0) := x"5DB26C4773E41517D7AABEB74D476462A5653E51F68C8B2F3A042766A18D0CA5";
   constant CPIX_NORMAL_INIT_72_BIT_09_C : bit_vector(255 downto 0) := x"12C1D4CF15149865E852D911C48CBAA445EDD862F9E8FF44FEDB6E4E151E0239";
   constant CPIX_NORMAL_INIT_72_BIT_10_C : bit_vector(255 downto 0) := x"C94C413FCDBFCF98CF32DA6F180C822C6C671BE7E57BC84FA3F58D5C3A5CB8C3";
   constant CPIX_NORMAL_INIT_72_BIT_11_C : bit_vector(255 downto 0) := x"87A5777C696629C7AE9C33667BF33B240ADC1D0ABE3B49A28B3FF026E5BC585F";
   constant CPIX_NORMAL_INIT_72_BIT_12_C : bit_vector(255 downto 0) := x"A90EAD356A9EF8486DB2A7256D855DFB664401E7EEC91DB9793FEE5D106E413D";
   constant CPIX_NORMAL_INIT_72_BIT_13_C : bit_vector(255 downto 0) := x"BBF43133276F5A2235F5EA0E241C4BF25CAE956188F2ADC10651B1ACE1559AFC";
   constant CPIX_NORMAL_INIT_72_BIT_14_C : bit_vector(255 downto 0) := x"234393B87DDCF3FE092A943D20A580C41634677E39FA0CFADE3D1390DB810F0A";
   constant CPIX_NORMAL_INIT_73_BIT_00_C : bit_vector(255 downto 0) := x"4016FD55357916D03A138450AD9C1E9F134CC5E31A4990A465B7CF08592A0C91";
   constant CPIX_NORMAL_INIT_73_BIT_01_C : bit_vector(255 downto 0) := x"15E62A0205450D725D3F151B41062BD566E7723D3D8C9A9B73B2381250452A61";
   constant CPIX_NORMAL_INIT_73_BIT_02_C : bit_vector(255 downto 0) := x"05347B52E13D34E4FB7313EC6D28D0D8688AC81689C795835502102025714672";
   constant CPIX_NORMAL_INIT_73_BIT_03_C : bit_vector(255 downto 0) := x"B0DA8643B0031F533A52A6856B235843D93DC11C26A5D5F91DC0A32B51321335";
   constant CPIX_NORMAL_INIT_73_BIT_04_C : bit_vector(255 downto 0) := x"574A331F504D29557B8AEF33F5BC60A68F7A7CCC4C9A35883B60A036915B5FA2";
   constant CPIX_NORMAL_INIT_73_BIT_05_C : bit_vector(255 downto 0) := x"D2714AA47CA495DA71D9D2B036766339DB191461247ABD2BEDEA9DE74EC7E01E";
   constant CPIX_NORMAL_INIT_73_BIT_06_C : bit_vector(255 downto 0) := x"1A051271E5455F7505A08D7B4A1244D7241D3A8E5A670EE8FE7CE55C920C1636";
   constant CPIX_NORMAL_INIT_73_BIT_07_C : bit_vector(255 downto 0) := x"175BD1678FDC41B01CE6E581FDCF4F33D4425A50668CB4946A5D4727C7702246";
   constant CPIX_NORMAL_INIT_73_BIT_08_C : bit_vector(255 downto 0) := x"49475270BC304F62A6B27AC177BCA2A7CA0BEF53BC23739B5C9D354B86160711";
   constant CPIX_NORMAL_INIT_73_BIT_09_C : bit_vector(255 downto 0) := x"0DB26359780DB36A391107CE835BD68A13F6CB2C12BD6199777B133EE4707701";
   constant CPIX_NORMAL_INIT_73_BIT_10_C : bit_vector(255 downto 0) := x"1CC67215093B06ACB50721C3A06C798D581FB231AB6C444430D2840E10172443";
   constant CPIX_NORMAL_INIT_73_BIT_11_C : bit_vector(255 downto 0) := x"7F933010C06C296B5210957982A583E260F3A509CBC0174C4E4206597044AAE8";
   constant CPIX_NORMAL_INIT_73_BIT_12_C : bit_vector(255 downto 0) := x"15C726248012359E72C973328A3C383AB76D526ECA1AE26804708724E9BA64BA";
   constant CPIX_NORMAL_INIT_73_BIT_13_C : bit_vector(255 downto 0) := x"52111644A7046ED4253FE1DC7D7A37537533CC98854C88C329D1BBBD7D0D6D7F";
   constant CPIX_NORMAL_INIT_73_BIT_14_C : bit_vector(255 downto 0) := x"4957E9CE9440173006D57DEC7F4A8EABE454AA191DB569717E32EB222F0D4969";
   constant CPIX_NORMAL_INIT_74_BIT_00_C : bit_vector(255 downto 0) := x"04A77C7FCA86855E375F9BD8414BDC1A561826669D1C6E098F624D99764BA343";
   constant CPIX_NORMAL_INIT_74_BIT_01_C : bit_vector(255 downto 0) := x"F23953F21509FBA49150D9D3699D4FE8F5A907A89372BB77FE1CD47DC4C52A29";
   constant CPIX_NORMAL_INIT_74_BIT_02_C : bit_vector(255 downto 0) := x"D11A3B5F09EBD2FA59A3ADCDE0425B33D1FB9B6F0B83C1FC04B06EB9455AB246";
   constant CPIX_NORMAL_INIT_74_BIT_03_C : bit_vector(255 downto 0) := x"4928A3B9AF09D4A17FA563A2F754D0226F77CF082263ECDBB8C7504B2F4A5A1F";
   constant CPIX_NORMAL_INIT_74_BIT_04_C : bit_vector(255 downto 0) := x"95AFF07518828647E7E948FCBD3387C7980E08675CCD5E2B7F48EE0BA5CA4499";
   constant CPIX_NORMAL_INIT_74_BIT_05_C : bit_vector(255 downto 0) := x"04CC5098A8A02043D5A4C7CF0F27EDB5231F347288182EA61B6EF05DF3CEE8C8";
   constant CPIX_NORMAL_INIT_74_BIT_06_C : bit_vector(255 downto 0) := x"2147A059AE62B8CA047700AE3D1A7ADC045F50F380F0C21A3FFBEF384EC46FAE";
   constant CPIX_NORMAL_INIT_74_BIT_07_C : bit_vector(255 downto 0) := x"0FFA48BA5AF0D87B623CBB3D6A703ECE2196A8D251B93F55FA82BC2736F9723F";
   constant CPIX_NORMAL_INIT_74_BIT_08_C : bit_vector(255 downto 0) := x"0D0BFC385606C654B8039656F306F4282A5D4413E0401D9BD1106240ED7FC9BF";
   constant CPIX_NORMAL_INIT_74_BIT_09_C : bit_vector(255 downto 0) := x"256C2872D7F8E31708BB57820057922D2C0AF88085CB00148FF789BCFB4490CB";
   constant CPIX_NORMAL_INIT_74_BIT_10_C : bit_vector(255 downto 0) := x"CEFB5EA69C19A2EB1355C927F063B963E2326569AA87EA7F27E56BB08653F78E";
   constant CPIX_NORMAL_INIT_74_BIT_11_C : bit_vector(255 downto 0) := x"602B912BC6F5C3D94FBCF623DFAB9E738C1FB73CC85372C1111F364D963E437C";
   constant CPIX_NORMAL_INIT_74_BIT_12_C : bit_vector(255 downto 0) := x"330048F33261209F7D825B40AD03F7ACF2E687B2B0BB7EEEFD031B1A135D13DC";
   constant CPIX_NORMAL_INIT_74_BIT_13_C : bit_vector(255 downto 0) := x"2D86B8802D92AF91026D15C81C9BEA5FDF0B4771570F3DE3D90719B0191DE4B7";
   constant CPIX_NORMAL_INIT_74_BIT_14_C : bit_vector(255 downto 0) := x"664EA79ECEB58C444D07711D7B0A726B7C563DA57D9532289881599B6AE3B780";
   constant CPIX_NORMAL_INIT_75_BIT_00_C : bit_vector(255 downto 0) := x"40D200BA0C2C5023EC66BBA8174692A00C234273304FB2C66D3659A18DA866A6";
   constant CPIX_NORMAL_INIT_75_BIT_01_C : bit_vector(255 downto 0) := x"F7A43DE1B895967F6389D7AF958A0BBFF8E1F6E9CB362D8D8230DE820770A5C3";
   constant CPIX_NORMAL_INIT_75_BIT_02_C : bit_vector(255 downto 0) := x"B7B36DD6B7EC2F5EDF40CD0E4BDF32B3BDC4E67AC272A88DD1DC08205BF90E1B";
   constant CPIX_NORMAL_INIT_75_BIT_03_C : bit_vector(255 downto 0) := x"6F586D4472EA978E076293DB56DE9C4729A4A7ADE03CC9790AB52CC93EF87198";
   constant CPIX_NORMAL_INIT_75_BIT_04_C : bit_vector(255 downto 0) := x"D49FB0E2CF6491C3B7E6EFC8C91BAE2B9E18F92301CA3226191ADD8555F79515";
   constant CPIX_NORMAL_INIT_75_BIT_05_C : bit_vector(255 downto 0) := x"A477497AEC9273ADE94D4DE60748DA70A1B766088D6E98136047255ADBD37B1D";
   constant CPIX_NORMAL_INIT_75_BIT_06_C : bit_vector(255 downto 0) := x"27840109934FB9065A79364771BFF20E870CA5E0E4B2E11197927C369D272E37";
   constant CPIX_NORMAL_INIT_75_BIT_07_C : bit_vector(255 downto 0) := x"6D76C38C8D20863ED76EDA7C6A5989188255E4016CA7D78C8174122E2E9915EA";
   constant CPIX_NORMAL_INIT_75_BIT_08_C : bit_vector(255 downto 0) := x"22C08164C50EB287DD9C3C3FDD4998B7C6248554712CE058CF76C6B76815F2C1";
   constant CPIX_NORMAL_INIT_75_BIT_09_C : bit_vector(255 downto 0) := x"4ACBB235F3D55B22F8CDE56453966C2C0214B1911E75610D2CCDA7C72C712C3F";
   constant CPIX_NORMAL_INIT_75_BIT_10_C : bit_vector(255 downto 0) := x"035C9234A96D63F12C13D9A3F9D6DC794031604478DAE4A802F015B596699625";
   constant CPIX_NORMAL_INIT_75_BIT_11_C : bit_vector(255 downto 0) := x"36580219637BA9B159EDCC9D2C9633C93BFF318027D2B064184F2698366DA71A";
   constant CPIX_NORMAL_INIT_75_BIT_12_C : bit_vector(255 downto 0) := x"405E0755EE71E1426753E6215C2CC37C7B11BB6B289785C4FD23F544A7BCCF70";
   constant CPIX_NORMAL_INIT_75_BIT_13_C : bit_vector(255 downto 0) := x"0480102D8E57F584C65D7AF759F7289973125A2012883FFE39D53A835CC2C8B6";
   constant CPIX_NORMAL_INIT_75_BIT_14_C : bit_vector(255 downto 0) := x"4344EE9A8545C9926DA756662D882D73370276363F41C396D90026B6973B6A8D";
   constant CPIX_NORMAL_INIT_76_BIT_00_C : bit_vector(255 downto 0) := x"0C0D817A677AF5084FFF50E7094B35805E5E4093744D91624A3AC41D3AE5B08F";
   constant CPIX_NORMAL_INIT_76_BIT_01_C : bit_vector(255 downto 0) := x"B174FCE8A9BDCE8346C3685FBAFFA63BEE6BB3445EE7AD7DE39B11EED378A37D";
   constant CPIX_NORMAL_INIT_76_BIT_02_C : bit_vector(255 downto 0) := x"9F707CDE8A4DBE478BD0E1615DDE07AAA4E8B95D7FBD6F2E0E281B0B94B261E1";
   constant CPIX_NORMAL_INIT_76_BIT_03_C : bit_vector(255 downto 0) := x"6B17BFA1391D13A787A1D79A22507D923046BC6F5BB72FAF09AFB6704D44A7CA";
   constant CPIX_NORMAL_INIT_76_BIT_04_C : bit_vector(255 downto 0) := x"DC07CF1844382CC8B28778C6EF11E42FD71608BEF0A823A2BADBBDE4381EE96E";
   constant CPIX_NORMAL_INIT_76_BIT_05_C : bit_vector(255 downto 0) := x"05A7C62FC502A8BCBAA3F898DD3AE8F9478D478DE19082B0A44C78C0DD7A7A08";
   constant CPIX_NORMAL_INIT_76_BIT_06_C : bit_vector(255 downto 0) := x"6C8ED7ADF18811602FBE9F6A5BCCB42E098DAB78302A8363307D08CB6A7B977F";
   constant CPIX_NORMAL_INIT_76_BIT_07_C : bit_vector(255 downto 0) := x"06E74760E7F0DABD7D332DD27B29FFA2492229C1B580066A0F2356AEF8AB107E";
   constant CPIX_NORMAL_INIT_76_BIT_08_C : bit_vector(255 downto 0) := x"867C23DD89ECD74A94E39AD4060BB3E8ABDCFE8C735B1C863D5B7FE04A2CEDAE";
   constant CPIX_NORMAL_INIT_76_BIT_09_C : bit_vector(255 downto 0) := x"42BE0E87FA57D4BA33C26C151FD759AF804335A3990CC64362514711AFFB840C";
   constant CPIX_NORMAL_INIT_76_BIT_10_C : bit_vector(255 downto 0) := x"023B88E0C1E6683A38C494CC92C6B619CA0C5AC68DD80680C7BDF0A70DE512BF";
   constant CPIX_NORMAL_INIT_76_BIT_11_C : bit_vector(255 downto 0) := x"489249A1115C799DC28C2E82E50D3AB08A811F2D2848BDBE400F8EB9628B9628";
   constant CPIX_NORMAL_INIT_76_BIT_12_C : bit_vector(255 downto 0) := x"4F038B2066FD95DE618B7277DBA22EEE4749462873BFC2BF08C451CBC6795FA1";
   constant CPIX_NORMAL_INIT_76_BIT_13_C : bit_vector(255 downto 0) := x"329D4165D362BD84C533E6D1B4892445377B4B8F5D5F730D5EBA49C2243DE6F8";
   constant CPIX_NORMAL_INIT_76_BIT_14_C : bit_vector(255 downto 0) := x"6F0C7E7F479AADF8F8255DA42C50668210D87710D417D35D3383AA7FBC8D4C7D";
   constant CPIX_NORMAL_INIT_77_BIT_00_C : bit_vector(255 downto 0) := x"455027AE2F06202C8294EF94D3023D88036815B317344DA279B2C750C62A0231";
   constant CPIX_NORMAL_INIT_77_BIT_01_C : bit_vector(255 downto 0) := x"D8F4F777ACB4B8DBAFAB4812D94B801CD2B6C266F6C4FCBC8C7E536BD75265F1";
   constant CPIX_NORMAL_INIT_77_BIT_02_C : bit_vector(255 downto 0) := x"315760273051644B439942EB0E7B57585E592D995675263EA2E331B5B8E84290";
   constant CPIX_NORMAL_INIT_77_BIT_03_C : bit_vector(255 downto 0) := x"E6CF51CC6D7D5E78592DB986EBA1007A0206587D61763D331B7879239485BFA8";
   constant CPIX_NORMAL_INIT_77_BIT_04_C : bit_vector(255 downto 0) := x"917D8987BDCAB9A9493360A061821F81B3A184B798ABC68AE83BEBD38D78D34D";
   constant CPIX_NORMAL_INIT_77_BIT_05_C : bit_vector(255 downto 0) := x"280713014F0B6E232229119BD8CFB67F452B0E1611334C4CBEF4232FBE17B2BE";
   constant CPIX_NORMAL_INIT_77_BIT_06_C : bit_vector(255 downto 0) := x"3931244433633F1A5C30EAC3D7398270BAFE77393F2E1748D04BF3D3F4D5A401";
   constant CPIX_NORMAL_INIT_77_BIT_07_C : bit_vector(255 downto 0) := x"2AF71B33004C9BE0B2D23973877598805DD21B370C35313FCAD0C55FF8468C57";
   constant CPIX_NORMAL_INIT_77_BIT_08_C : bit_vector(255 downto 0) := x"457330075B4A3C8C6F9D8A583966ED5C72E41D6C1F016F18663CBD694B66C8D7";
   constant CPIX_NORMAL_INIT_77_BIT_09_C : bit_vector(255 downto 0) := x"425D352BB8DE1B8A9CF3DC431E8275FD7FEF3B607A60254339ADF47BDCC83B60";
   constant CPIX_NORMAL_INIT_77_BIT_10_C : bit_vector(255 downto 0) := x"6717321A5B8820A4C49A83AF04231A3861030F4547276B01C9CA0642BD6D7E97";
   constant CPIX_NORMAL_INIT_77_BIT_11_C : bit_vector(255 downto 0) := x"6A30240D45FF07079929CD71B6BE35570B43315189DA475ECC12476592A0BC5F";
   constant CPIX_NORMAL_INIT_77_BIT_12_C : bit_vector(255 downto 0) := x"2267031966806950CCDD69C93C4CC54E024F162502CCADBF9DC0111A399F537D";
   constant CPIX_NORMAL_INIT_77_BIT_13_C : bit_vector(255 downto 0) := x"297152454B46422867CA6C2CC0C27E6C4166B2B856FE46BEC386D8C596D1683E";
   constant CPIX_NORMAL_INIT_77_BIT_14_C : bit_vector(255 downto 0) := x"0077CBAF3A0805047AC28DD1338BF7542B0C4CFA04EA07FD362874AEC9E4670F";
   constant CPIX_NORMAL_INIT_78_BIT_00_C : bit_vector(255 downto 0) := x"E39B2798F279B802D5AE3365A2DBFB86D41BEDAB45BF4E105F20A7DACFEDC5BA";
   constant CPIX_NORMAL_INIT_78_BIT_01_C : bit_vector(255 downto 0) := x"DFEF6CB9E2E44A5C86E563DF2A7AE552C9D5C8C74B87DE971EB6D008A2F8CD9C";
   constant CPIX_NORMAL_INIT_78_BIT_02_C : bit_vector(255 downto 0) := x"F3FB655E54A6826D123C8BE02B3BCDAB5FEE28417B8167CA8CE8714D55213437";
   constant CPIX_NORMAL_INIT_78_BIT_03_C : bit_vector(255 downto 0) := x"248EF65E28EFFD042642BD1D32BADF320059446754CE466C6EBF03AF1F4B4BF3";
   constant CPIX_NORMAL_INIT_78_BIT_04_C : bit_vector(255 downto 0) := x"2BB2E6BE4ACCBECD1A617485715DF58A390F5547E4EA5A94F97C835826717BAB";
   constant CPIX_NORMAL_INIT_78_BIT_05_C : bit_vector(255 downto 0) := x"3D836C9B900776E78BEA1CE8B199C91F07775C239018744ED7987CE11A5A1F91";
   constant CPIX_NORMAL_INIT_78_BIT_06_C : bit_vector(255 downto 0) := x"3117271D6936CDBB4DC8EBEB7B3D6A96EA403D3DD50AB52583B3A305653E0ACF";
   constant CPIX_NORMAL_INIT_78_BIT_07_C : bit_vector(255 downto 0) := x"1607CADF6EAB156E36F14B2BE139452F517C4A59C1708DCD607EC054099C6C7B";
   constant CPIX_NORMAL_INIT_78_BIT_08_C : bit_vector(255 downto 0) := x"BBD4F9843C86E5A05DCF9A194CA1B8DC631C380D23F9DF573C58993E698A4C64";
   constant CPIX_NORMAL_INIT_78_BIT_09_C : bit_vector(255 downto 0) := x"2AB8DA7B75BD10A6250598EEC82056207F0E150AD90EDF9AD7395FA8C9AC5651";
   constant CPIX_NORMAL_INIT_78_BIT_10_C : bit_vector(255 downto 0) := x"2E880AB5E142D99ABEB36E9C99806119041C2435DFFB31AD98A46A2068926877";
   constant CPIX_NORMAL_INIT_78_BIT_11_C : bit_vector(255 downto 0) := x"008D4C549CCA30910CC8FAA309FE7E88254639ECE27A3769CE4D55F21F341C4B";
   constant CPIX_NORMAL_INIT_78_BIT_12_C : bit_vector(255 downto 0) := x"340CD9D3E2BA67A701A576416EF13A052D109E904C55488C9D8F991A304F2C32";
   constant CPIX_NORMAL_INIT_78_BIT_13_C : bit_vector(255 downto 0) := x"6C15D025DC12B5657AADBB525D172C6603C23AF1F57BC5B5391B7BA12101654E";
   constant CPIX_NORMAL_INIT_78_BIT_14_C : bit_vector(255 downto 0) := x"387B9BE511A3521B647A1F9AD45570C028E93FA083375A0261CCF1A66814AE70";
   constant CPIX_NORMAL_INIT_79_BIT_00_C : bit_vector(255 downto 0) := x"FE1FB9E78E7F15C4ED72CD73B24DD8D787CDC3A382D9E3D3823327DA5F8BA04F";
   constant CPIX_NORMAL_INIT_79_BIT_01_C : bit_vector(255 downto 0) := x"F36EB9C2A97C14BCB024A7C8EF2CD8A3A6B6DB38E82CC377BC21E3FAFCEB3CF3";
   constant CPIX_NORMAL_INIT_79_BIT_02_C : bit_vector(255 downto 0) := x"F67F7F8E7D62720ECB812CC9A3089C96973CAFE80C3022C807527E260FF52E65";
   constant CPIX_NORMAL_INIT_79_BIT_03_C : bit_vector(255 downto 0) := x"399FF8B379B86525268258CE8ADF9D967F0D9D26287B51BA362BC256BC81EF0D";
   constant CPIX_NORMAL_INIT_79_BIT_04_C : bit_vector(255 downto 0) := x"235D3AE273D5CE49B76A2B0AF6CD1BBF37C78166773E4FF000A24A90BFCF384B";
   constant CPIX_NORMAL_INIT_79_BIT_05_C : bit_vector(255 downto 0) := x"B43054094A9C5556B20447E76DA521411BA5B32E8FB58ECCD297DCAC3DED70DB";
   constant CPIX_NORMAL_INIT_79_BIT_06_C : bit_vector(255 downto 0) := x"1014D0340CA73109427B353EF6C292150E6429E6378BB82E17B221EE8E67BD7D";
   constant CPIX_NORMAL_INIT_79_BIT_07_C : bit_vector(255 downto 0) := x"1385AA0C2DC8EB3581305AC87215945102EE74E37973D6AB2A5C79CB6F2C3AA5";
   constant CPIX_NORMAL_INIT_79_BIT_08_C : bit_vector(255 downto 0) := x"2114E435DD785EDDB3F1E55B2A4391102F655C219FFD2145C470DAB77C55EA2D";
   constant CPIX_NORMAL_INIT_79_BIT_09_C : bit_vector(255 downto 0) := x"2D5262D7601B939B1DB61E4A5717C4501A8F0084E1A08AFC0EA5EEF0F7732317";
   constant CPIX_NORMAL_INIT_79_BIT_10_C : bit_vector(255 downto 0) := x"2950271EC149C66A23D4F60049830141A003AFBAB5B72296653DC7A3D8A252E8";
   constant CPIX_NORMAL_INIT_79_BIT_11_C : bit_vector(255 downto 0) := x"7940866710869C9D4DC2B812311240FE9C566569FA557D743A23F72DB7C5CE23";
   constant CPIX_NORMAL_INIT_79_BIT_12_C : bit_vector(255 downto 0) := x"0954814B5A55B667D617B3D60494EF4FE3E47BE26DD4682F500DFA2E67F20706";
   constant CPIX_NORMAL_INIT_79_BIT_13_C : bit_vector(255 downto 0) := x"1010D07847CA675145AA82A968FE6267FC4557354CF3423D2F84ADE810CEC0BE";
   constant CPIX_NORMAL_INIT_79_BIT_14_C : bit_vector(255 downto 0) := x"21EB8014186E73BFC0F22C6475F57226519E6ADF27864C8814576F2FB618B833";
   constant CPIX_NORMAL_INIT_7A_BIT_00_C : bit_vector(255 downto 0) := x"F6F0D9FA1A01EE63DAEABC269AD351A2F298467CAC45FC5CEDAA5D8D4AD5AC2E";
   constant CPIX_NORMAL_INIT_7A_BIT_01_C : bit_vector(255 downto 0) := x"2A9C316D409E655C3634094C0E6A456B248544802CEC966223B4C878B8532458";
   constant CPIX_NORMAL_INIT_7A_BIT_02_C : bit_vector(255 downto 0) := x"FFF9CF1BB0A35F1DFAF79DEE80667F11A3F36B9F01AE5575AE177186042F27D9";
   constant CPIX_NORMAL_INIT_7A_BIT_03_C : bit_vector(255 downto 0) := x"50F05E93159B5FA17EFECEA23C283F4A065EB28C7C59C4C555B215EBE902573B";
   constant CPIX_NORMAL_INIT_7A_BIT_04_C : bit_vector(255 downto 0) := x"8B5DB489DDFAE7F7A0C5035523A80C808FC42991DE2EE1D9A3252A3772F3CF02";
   constant CPIX_NORMAL_INIT_7A_BIT_05_C : bit_vector(255 downto 0) := x"C537E95EE22D56B4CD52A7A14143B9720A0AEC418C9B35AC5345A27D37C2DFEA";
   constant CPIX_NORMAL_INIT_7A_BIT_06_C : bit_vector(255 downto 0) := x"581293E136510BD392CCCDC09965A57541C2F5EB050F637A030D8C937FF63C7F";
   constant CPIX_NORMAL_INIT_7A_BIT_07_C : bit_vector(255 downto 0) := x"658AA49797B672A290C06D9A84177A0F3F2F3CA756F6747B49E90E70F9E55A57";
   constant CPIX_NORMAL_INIT_7A_BIT_08_C : bit_vector(255 downto 0) := x"588483D9AA67A2AD948046C2B59D60D823E61190E191D1C67201C02B8050E7AF";
   constant CPIX_NORMAL_INIT_7A_BIT_09_C : bit_vector(255 downto 0) := x"3BD4D835EAC4196610C834426AD9646746659ED12F19019663E88B00BDAEF08B";
   constant CPIX_NORMAL_INIT_7A_BIT_10_C : bit_vector(255 downto 0) := x"1294E65C61ADE9A604406BCE1C0C9694BF3DA2DF10A5C5E5D546F9F75C7C91DB";
   constant CPIX_NORMAL_INIT_7A_BIT_11_C : bit_vector(255 downto 0) := x"521257EC2EAA695A7F4859C4235A56D347879C9A3ED5BFB5A3D6A15803529716";
   constant CPIX_NORMAL_INIT_7A_BIT_12_C : bit_vector(255 downto 0) := x"0310F4C151D4269670F76988E5C0DEB4502D544B6930E1DEDD9DCF7FE133121A";
   constant CPIX_NORMAL_INIT_7A_BIT_13_C : bit_vector(255 downto 0) := x"0806B1C8927D2D6A51341A7F687929AD69E869F8160A2BF3B314136DA12C22CD";
   constant CPIX_NORMAL_INIT_7A_BIT_14_C : bit_vector(255 downto 0) := x"10FB80A96D156A6551557099A05D977A53DBBCA021427357616C6856A82B7DD8";
   constant CPIX_NORMAL_INIT_7B_BIT_00_C : bit_vector(255 downto 0) := x"FFA08EB967076E95E9F2EBD2926F68EBDD78A83DC0F2DCB7CCF6BD7AC87D8334";
   constant CPIX_NORMAL_INIT_7B_BIT_01_C : bit_vector(255 downto 0) := x"537562529826CD177467333C3578F9A719964684D99123603B26809C137215E2";
   constant CPIX_NORMAL_INIT_7B_BIT_02_C : bit_vector(255 downto 0) := x"126542531A197B0752083747CD2486BBAD7BB2F578542B3FC6C4FE6F36438C6C";
   constant CPIX_NORMAL_INIT_7B_BIT_03_C : bit_vector(255 downto 0) := x"C92A642626E9B402512666653645885D78EC6219DC8B504941E3BD772F9420FB";
   constant CPIX_NORMAL_INIT_7B_BIT_04_C : bit_vector(255 downto 0) := x"8689EBEE254C49389C8D8D9BE7F9A693A9B2066A9969F0C7912F4E5DFBEC63C7";
   constant CPIX_NORMAL_INIT_7B_BIT_05_C : bit_vector(255 downto 0) := x"61103375560BABD707310522FC57F1DE059781EEFDEAA7EE1A1AC89CC268A772";
   constant CPIX_NORMAL_INIT_7B_BIT_06_C : bit_vector(255 downto 0) := x"6440557324F99694FF56771283D9C8C06B9ECA047FB73AC72AF64795462B7797";
   constant CPIX_NORMAL_INIT_7B_BIT_07_C : bit_vector(255 downto 0) := x"7D3502BCD96594A829352447B883E1A11D14DCBE656976FD2568C817351FEF07";
   constant CPIX_NORMAL_INIT_7B_BIT_08_C : bit_vector(255 downto 0) := x"0541336A7AB265E25C26307256E635A9965AAE938DB813DEFAFA5329637C36EF";
   constant CPIX_NORMAL_INIT_7B_BIT_09_C : bit_vector(255 downto 0) := x"1247EB3BADA1394E7F7474416EC7AA741F39F18F5960392F814DA2915010FF82";
   constant CPIX_NORMAL_INIT_7B_BIT_10_C : bit_vector(255 downto 0) := x"51533A4C8B9F053641301570AB11E67917AC8D67688A99D2B239AA189ECD2C1F";
   constant CPIX_NORMAL_INIT_7B_BIT_11_C : bit_vector(255 downto 0) := x"74420F11A6A4DF413140AB13A1149CE3292C026A9A79C27CB83662EF03BE5B96";
   constant CPIX_NORMAL_INIT_7B_BIT_12_C : bit_vector(255 downto 0) := x"55125860AA6A628313141AEFA8036B1631B45E8B4B55BD7F12165F9F280B963C";
   constant CPIX_NORMAL_INIT_7B_BIT_13_C : bit_vector(255 downto 0) := x"641031165B66897605DE1F1F99A898675A0495E885D8CA40573B23523F2946DE";
   constant CPIX_NORMAL_INIT_7B_BIT_14_C : bit_vector(255 downto 0) := x"05BF720079A85BD0722F0F1E564FAC5372771BEEE42C60590A50819259F7EA26";
   constant CPIX_NORMAL_INIT_7C_BIT_00_C : bit_vector(255 downto 0) := x"0C1248F71A5A2D56656265266AA4C43C24A5291E70AB24067C10F0CFCB244170";
   constant CPIX_NORMAL_INIT_7C_BIT_01_C : bit_vector(255 downto 0) := x"DBFBAEF9DE80DBFBB8D483B38E7B2B519BCBF52CECF053C7D4B9C976F6A69FDA";
   constant CPIX_NORMAL_INIT_7C_BIT_02_C : bit_vector(255 downto 0) := x"DF696DA2A26ADBFBB6BE25781B553C64DFC22C9A761C77A96B70B81D6C660515";
   constant CPIX_NORMAL_INIT_7C_BIT_03_C : bit_vector(255 downto 0) := x"63ED66E45B2BB2FB52A5662F5D91E8F24B534FE831E25FB542158B123F3B322D";
   constant CPIX_NORMAL_INIT_7C_BIT_04_C : bit_vector(255 downto 0) := x"527D5812D573DA6D5985571C0538FB637DDF3AF2144842CB23114F38E6B2547F";
   constant CPIX_NORMAL_INIT_7C_BIT_05_C : bit_vector(255 downto 0) := x"C4023A01D01D6C003CD7BCBA99AE6E4B696B815DBF2ECAA3153582439A4C3338";
   constant CPIX_NORMAL_INIT_7C_BIT_06_C : bit_vector(255 downto 0) := x"00842D421747D990346D5BE71D4FB5E6415265AF2AFF7679F07683C49DD0473B";
   constant CPIX_NORMAL_INIT_7C_BIT_07_C : bit_vector(255 downto 0) := x"18F26AF4843A50801F4D659F726B767C11BB7F075C37C607062284AA47802A67";
   constant CPIX_NORMAL_INIT_7C_BIT_08_C : bit_vector(255 downto 0) := x"40C4A63ADCC371807424BE4084BD60F6F8E869CC2BB22CEA52625EB162A76B24";
   constant CPIX_NORMAL_INIT_7C_BIT_09_C : bit_vector(255 downto 0) := x"6159439B2D3311803B08CCBE3CFCD5517EB74E0D40AFA4147303A3BB963EAE10";
   constant CPIX_NORMAL_INIT_7C_BIT_10_C : bit_vector(255 downto 0) := x"6053829758D02900C1FFCD59469DAD1E7A3CC1ABFD7AA8420244BF4EAC746965";
   constant CPIX_NORMAL_INIT_7C_BIT_11_C : bit_vector(255 downto 0) := x"609509AA29E1410FA146F06475D6D8B50A20AB482AFD2F7A416ED756B20D3423";
   constant CPIX_NORMAL_INIT_7C_BIT_12_C : bit_vector(255 downto 0) := x"208330D591D908F3DC7D686702F75D1142A9DF5D0C507C7060B8202AABA34365";
   constant CPIX_NORMAL_INIT_7C_BIT_13_C : bit_vector(255 downto 0) := x"00861B500F9E6F55E0142D1678EE0B8F6084A1C47EF12165197CC78C637C4043";
   constant CPIX_NORMAL_INIT_7C_BIT_14_C : bit_vector(255 downto 0) := x"4F80275F8D644C550B7B592A0177D2E567BC0D13473B80486E7C95314ACD60F4";
   constant CPIX_NORMAL_INIT_7D_BIT_00_C : bit_vector(255 downto 0) := x"0341AE8712066890591972525218596B2350CF0A401A46F225E91F1D10D5C718";
   constant CPIX_NORMAL_INIT_7D_BIT_01_C : bit_vector(255 downto 0) := x"17100B2657502E7D7001DA0627924C665916C448143871F56DE171884C73265A";
   constant CPIX_NORMAL_INIT_7D_BIT_02_C : bit_vector(255 downto 0) := x"1711387700518C8FB7DD32759AE719C4FFA3093AFDB7C580F89A1E0CF1180142";
   constant CPIX_NORMAL_INIT_7D_BIT_03_C : bit_vector(255 downto 0) := x"A44556C7055458A27E53B9020FE5700F0D390B347FAD26F3335A72800D1FE117";
   constant CPIX_NORMAL_INIT_7D_BIT_04_C : bit_vector(255 downto 0) := x"9AFF4220AAABD6D9FD16B6C98532FE59B3CAAFDDC8105EA89868A7CAD4655DB1";
   constant CPIX_NORMAL_INIT_7D_BIT_05_C : bit_vector(255 downto 0) := x"405413F91405E1CB198FFFDF33AA96D584E3D61CA1DC016533E0AB4E10D659BF";
   constant CPIX_NORMAL_INIT_7D_BIT_06_C : bit_vector(255 downto 0) := x"40054E98F1519AA86BB06D797D181759219C50399AA8A4C409CF035712A97D67";
   constant CPIX_NORMAL_INIT_7D_BIT_07_C : bit_vector(255 downto 0) := x"641EA48E6441E9CC20AF465E46A143F14BC99D5D886B8173776D1D472E34EC31";
   constant CPIX_NORMAL_INIT_7D_BIT_08_C : bit_vector(255 downto 0) := x"00577D4D25451D4E93F9AE1BFF16565F289AF5DE8819CA4A5D08C889508780DF";
   constant CPIX_NORMAL_INIT_7D_BIT_09_C : bit_vector(255 downto 0) := x"11F7EC63744079F436CB246782D800F978A4F8250A417A4514B872095EB0EFCB";
   constant CPIX_NORMAL_INIT_7D_BIT_10_C : bit_vector(255 downto 0) := x"0172BB050404F0D61EA56BA9D6F2BA6318D24EED007B2298F6DB0C8C81ED268B";
   constant CPIX_NORMAL_INIT_7D_BIT_11_C : bit_vector(255 downto 0) := x"4130DCB040F1C0AD6617B696E55F1F39111E7F637228531919AB78FCD9C21191";
   constant CPIX_NORMAL_INIT_7D_BIT_12_C : bit_vector(255 downto 0) := x"0124F759103FE1714C3B30E7113B639610C808594D6AC8BC060364CBAAB7C513";
   constant CPIX_NORMAL_INIT_7D_BIT_13_C : bit_vector(255 downto 0) := x"404135A50B33AEA5308E8AB01751761B21CA96670437666E6E6E137DD016C65A";
   constant CPIX_NORMAL_INIT_7D_BIT_14_C : bit_vector(255 downto 0) := x"0F506E38573313E1553FC64230892DF50F8E6074004AC2971BEC41514661E76A";
   constant CPIX_NORMAL_INIT_7E_BIT_00_C : bit_vector(255 downto 0) := x"EF06EE97DDAEEDD8AF4CFCE2B1CDF76DDED2CC9EBABA8379B39CB0BE9F344BFB";
   constant CPIX_NORMAL_INIT_7E_BIT_01_C : bit_vector(255 downto 0) := x"FF33FEE19D1FB4FD8ECEFAAEDD87D23E612C742152273409085A5CA711919640";
   constant CPIX_NORMAL_INIT_7E_BIT_02_C : bit_vector(255 downto 0) := x"FF67EE2A475A19F0736B152A7AB7102DF66D93BFCD64306DB97342F865F26740";
   constant CPIX_NORMAL_INIT_7E_BIT_03_C : bit_vector(255 downto 0) := x"2F1BEE2D74EB3C93247C6E7F43DD33ED1E5C37DF1C7728E4312E4D9C11A17516";
   constant CPIX_NORMAL_INIT_7E_BIT_04_C : bit_vector(255 downto 0) := x"9016119AE5D08562DBB2A01CA65E9400162185B6283206F56B7D029B5136DD07";
   constant CPIX_NORMAL_INIT_7E_BIT_05_C : bit_vector(255 downto 0) := x"001C00CB2FFB5F988D92CA045CF7192F8170826069CFAF736782F73D0591B256";
   constant CPIX_NORMAL_INIT_7E_BIT_06_C : bit_vector(255 downto 0) := x"003AC0BE786662124A06BEC82B150E65086111A8463D23CD014F7F56C498A817";
   constant CPIX_NORMAL_INIT_7E_BIT_07_C : bit_vector(255 downto 0) := x"43CB40EA4F131C1C3AA2A785562574E42D7C8708324B57560F712591158F1875";
   constant CPIX_NORMAL_INIT_7E_BIT_08_C : bit_vector(255 downto 0) := x"016240239EF3F1136BCBA2B322AE098B08D7A94844F08E4DEE6A7D6F153C5D74";
   constant CPIX_NORMAL_INIT_7E_BIT_09_C : bit_vector(255 downto 0) := x"0DE5406C5B459A0E6CE430700E563CFB421B650872AF6E807D320FC051DF97F0";
   constant CPIX_NORMAL_INIT_7E_BIT_10_C : bit_vector(255 downto 0) := x"05F000C93C7E9DF5293E075ADB2E8E5B419928608FA21AE3768FE7E110F3E464";
   constant CPIX_NORMAL_INIT_7E_BIT_11_C : bit_vector(255 downto 0) := x"04AC0C8E51D9C336037556122F6AA908482F6C03C1C449AC34F27E770791D245";
   constant CPIX_NORMAL_INIT_7E_BIT_12_C : bit_vector(255 downto 0) := x"04D207C4274D07590A2227AE114BFD8149488A2DA6651D201EB220644E47FD14";
   constant CPIX_NORMAL_INIT_7E_BIT_13_C : bit_vector(255 downto 0) := x"004C35FC4BBC10534B9505577716819309303B70C0616F3B48C87C44269A5601";
   constant CPIX_NORMAL_INIT_7E_BIT_14_C : bit_vector(255 downto 0) := x"3076151C07914A6C3B4403993E0014D73853A4203727059C5E21178276843A4C";
   constant CPIX_NORMAL_INIT_7F_BIT_00_C : bit_vector(255 downto 0) := x"4F00FFFE40410106CEFFDEB9EFF9BBC70E0650150D1235294654006925304BC0";
   constant CPIX_NORMAL_INIT_7F_BIT_01_C : bit_vector(255 downto 0) := x"53F0FF010440FEEF31240016EFFEA9D7FBFAF3DBB6ED9CBE0010152B061D4350";
   constant CPIX_NORMAL_INIT_7F_BIT_02_C : bit_vector(255 downto 0) := x"57713F17E545477BFC321177743F6AF7FFF5433D5307692ED68FA46FE10E0E10";
   constant CPIX_NORMAL_INIT_7F_BIT_03_C : bit_vector(255 downto 0) := x"57717F176144567F6D16152537783FF779F60F7846771A76325B2545472A0E41";
   constant CPIX_NORMAL_INIT_7F_BIT_04_C : bit_vector(255 downto 0) := x"3B818056DEAA7779A3A8E99C2E7A7BDB890BC895BDC2D3A0148D651D761B07A1";
   constant CPIX_NORMAL_INIT_7F_BIT_05_C : bit_vector(255 downto 0) := x"05290CC355E4E00F3377EC61AC4401FB0A0B7F2AA9B02D0784946BF459D60AD1";
   constant CPIX_NORMAL_INIT_7F_BIT_06_C : bit_vector(255 downto 0) := x"01004401703051073B404F446713146F0F8F655131FA7034240E165A037188E1";
   constant CPIX_NORMAL_INIT_7F_BIT_07_C : bit_vector(255 downto 0) := x"010004401071601513456A027D104277130F31227DD8144C6692531134480B24";
   constant CPIX_NORMAL_INIT_7F_BIT_08_C : bit_vector(255 downto 0) := x"004234580E75268100E87A37492DD5570505BDC17BDD5F2B29E20CB2F7670624";
   constant CPIX_NORMAL_INIT_7F_BIT_09_C : bit_vector(255 downto 0) := x"0000100142410516614D6047113646792C0630B36C44316F13425F7865380B9C";
   constant CPIX_NORMAL_INIT_7F_BIT_10_C : bit_vector(255 downto 0) := x"00141325530A4D76235E51DD34E63A690C0A67AC6713B7B30A64BD3D5BDC0DC4";
   constant CPIX_NORMAL_INIT_7F_BIT_11_C : bit_vector(255 downto 0) := x"0004112156020D463738005D54A724690E2B0A95141177E22761882E4D751890";
   constant CPIX_NORMAL_INIT_7F_BIT_12_C : bit_vector(255 downto 0) := x"00040161501328422211431E5D84600D09185212355F03E822B6D4243D4431E0";
   constant CPIX_NORMAL_INIT_7F_BIT_13_C : bit_vector(255 downto 0) := x"00040120144308441370600A44857431024E3E0138015189247484772A605B10";
   constant CPIX_NORMAL_INIT_7F_BIT_14_C : bit_vector(255 downto 0) := x"0000004004112114012543424803422445021836701A700961C4550A34195872";

      
   
   
   
   
   
   
   
   
   
   
   type Bit256Array is array (natural range <>) of bit_vector(255 downto 0);
   
   
   constant CPIX_NORMAL_INIT_00_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_00_BIT_00_C, 1  => CPIX_NORMAL_INIT_00_BIT_01_C, 2  => CPIX_NORMAL_INIT_00_BIT_02_C, 3  => CPIX_NORMAL_INIT_00_BIT_03_C, 4  => CPIX_NORMAL_INIT_00_BIT_04_C, 5  => CPIX_NORMAL_INIT_00_BIT_05_C, 6  => CPIX_NORMAL_INIT_00_BIT_06_C, 7  => CPIX_NORMAL_INIT_00_BIT_07_C, 8  => CPIX_NORMAL_INIT_00_BIT_08_C, 9  => CPIX_NORMAL_INIT_00_BIT_09_C, 10 => CPIX_NORMAL_INIT_00_BIT_10_C, 11 => CPIX_NORMAL_INIT_00_BIT_11_C, 12 => CPIX_NORMAL_INIT_00_BIT_12_C, 13 => CPIX_NORMAL_INIT_00_BIT_13_C, 14 => CPIX_NORMAL_INIT_00_BIT_14_C);
   constant CPIX_NORMAL_INIT_01_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_01_BIT_00_C, 1  => CPIX_NORMAL_INIT_01_BIT_01_C, 2  => CPIX_NORMAL_INIT_01_BIT_02_C, 3  => CPIX_NORMAL_INIT_01_BIT_03_C, 4  => CPIX_NORMAL_INIT_01_BIT_04_C, 5  => CPIX_NORMAL_INIT_01_BIT_05_C, 6  => CPIX_NORMAL_INIT_01_BIT_06_C, 7  => CPIX_NORMAL_INIT_01_BIT_07_C, 8  => CPIX_NORMAL_INIT_01_BIT_08_C, 9  => CPIX_NORMAL_INIT_01_BIT_09_C, 10 => CPIX_NORMAL_INIT_01_BIT_10_C, 11 => CPIX_NORMAL_INIT_01_BIT_11_C, 12 => CPIX_NORMAL_INIT_01_BIT_12_C, 13 => CPIX_NORMAL_INIT_01_BIT_13_C, 14 => CPIX_NORMAL_INIT_01_BIT_14_C);
   constant CPIX_NORMAL_INIT_02_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_02_BIT_00_C, 1  => CPIX_NORMAL_INIT_02_BIT_01_C, 2  => CPIX_NORMAL_INIT_02_BIT_02_C, 3  => CPIX_NORMAL_INIT_02_BIT_03_C, 4  => CPIX_NORMAL_INIT_02_BIT_04_C, 5  => CPIX_NORMAL_INIT_02_BIT_05_C, 6  => CPIX_NORMAL_INIT_02_BIT_06_C, 7  => CPIX_NORMAL_INIT_02_BIT_07_C, 8  => CPIX_NORMAL_INIT_02_BIT_08_C, 9  => CPIX_NORMAL_INIT_02_BIT_09_C, 10 => CPIX_NORMAL_INIT_02_BIT_10_C, 11 => CPIX_NORMAL_INIT_02_BIT_11_C, 12 => CPIX_NORMAL_INIT_02_BIT_12_C, 13 => CPIX_NORMAL_INIT_02_BIT_13_C, 14 => CPIX_NORMAL_INIT_02_BIT_14_C);
   constant CPIX_NORMAL_INIT_03_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_03_BIT_00_C, 1  => CPIX_NORMAL_INIT_03_BIT_01_C, 2  => CPIX_NORMAL_INIT_03_BIT_02_C, 3  => CPIX_NORMAL_INIT_03_BIT_03_C, 4  => CPIX_NORMAL_INIT_03_BIT_04_C, 5  => CPIX_NORMAL_INIT_03_BIT_05_C, 6  => CPIX_NORMAL_INIT_03_BIT_06_C, 7  => CPIX_NORMAL_INIT_03_BIT_07_C, 8  => CPIX_NORMAL_INIT_03_BIT_08_C, 9  => CPIX_NORMAL_INIT_03_BIT_09_C, 10 => CPIX_NORMAL_INIT_03_BIT_10_C, 11 => CPIX_NORMAL_INIT_03_BIT_11_C, 12 => CPIX_NORMAL_INIT_03_BIT_12_C, 13 => CPIX_NORMAL_INIT_03_BIT_13_C, 14 => CPIX_NORMAL_INIT_03_BIT_14_C);
   constant CPIX_NORMAL_INIT_04_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_04_BIT_00_C, 1  => CPIX_NORMAL_INIT_04_BIT_01_C, 2  => CPIX_NORMAL_INIT_04_BIT_02_C, 3  => CPIX_NORMAL_INIT_04_BIT_03_C, 4  => CPIX_NORMAL_INIT_04_BIT_04_C, 5  => CPIX_NORMAL_INIT_04_BIT_05_C, 6  => CPIX_NORMAL_INIT_04_BIT_06_C, 7  => CPIX_NORMAL_INIT_04_BIT_07_C, 8  => CPIX_NORMAL_INIT_04_BIT_08_C, 9  => CPIX_NORMAL_INIT_04_BIT_09_C, 10 => CPIX_NORMAL_INIT_04_BIT_10_C, 11 => CPIX_NORMAL_INIT_04_BIT_11_C, 12 => CPIX_NORMAL_INIT_04_BIT_12_C, 13 => CPIX_NORMAL_INIT_04_BIT_13_C, 14 => CPIX_NORMAL_INIT_04_BIT_14_C);
   constant CPIX_NORMAL_INIT_05_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_05_BIT_00_C, 1  => CPIX_NORMAL_INIT_05_BIT_01_C, 2  => CPIX_NORMAL_INIT_05_BIT_02_C, 3  => CPIX_NORMAL_INIT_05_BIT_03_C, 4  => CPIX_NORMAL_INIT_05_BIT_04_C, 5  => CPIX_NORMAL_INIT_05_BIT_05_C, 6  => CPIX_NORMAL_INIT_05_BIT_06_C, 7  => CPIX_NORMAL_INIT_05_BIT_07_C, 8  => CPIX_NORMAL_INIT_05_BIT_08_C, 9  => CPIX_NORMAL_INIT_05_BIT_09_C, 10 => CPIX_NORMAL_INIT_05_BIT_10_C, 11 => CPIX_NORMAL_INIT_05_BIT_11_C, 12 => CPIX_NORMAL_INIT_05_BIT_12_C, 13 => CPIX_NORMAL_INIT_05_BIT_13_C, 14 => CPIX_NORMAL_INIT_05_BIT_14_C);
   constant CPIX_NORMAL_INIT_06_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_06_BIT_00_C, 1  => CPIX_NORMAL_INIT_06_BIT_01_C, 2  => CPIX_NORMAL_INIT_06_BIT_02_C, 3  => CPIX_NORMAL_INIT_06_BIT_03_C, 4  => CPIX_NORMAL_INIT_06_BIT_04_C, 5  => CPIX_NORMAL_INIT_06_BIT_05_C, 6  => CPIX_NORMAL_INIT_06_BIT_06_C, 7  => CPIX_NORMAL_INIT_06_BIT_07_C, 8  => CPIX_NORMAL_INIT_06_BIT_08_C, 9  => CPIX_NORMAL_INIT_06_BIT_09_C, 10 => CPIX_NORMAL_INIT_06_BIT_10_C, 11 => CPIX_NORMAL_INIT_06_BIT_11_C, 12 => CPIX_NORMAL_INIT_06_BIT_12_C, 13 => CPIX_NORMAL_INIT_06_BIT_13_C, 14 => CPIX_NORMAL_INIT_06_BIT_14_C);
   constant CPIX_NORMAL_INIT_07_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_07_BIT_00_C, 1  => CPIX_NORMAL_INIT_07_BIT_01_C, 2  => CPIX_NORMAL_INIT_07_BIT_02_C, 3  => CPIX_NORMAL_INIT_07_BIT_03_C, 4  => CPIX_NORMAL_INIT_07_BIT_04_C, 5  => CPIX_NORMAL_INIT_07_BIT_05_C, 6  => CPIX_NORMAL_INIT_07_BIT_06_C, 7  => CPIX_NORMAL_INIT_07_BIT_07_C, 8  => CPIX_NORMAL_INIT_07_BIT_08_C, 9  => CPIX_NORMAL_INIT_07_BIT_09_C, 10 => CPIX_NORMAL_INIT_07_BIT_10_C, 11 => CPIX_NORMAL_INIT_07_BIT_11_C, 12 => CPIX_NORMAL_INIT_07_BIT_12_C, 13 => CPIX_NORMAL_INIT_07_BIT_13_C, 14 => CPIX_NORMAL_INIT_07_BIT_14_C);
   constant CPIX_NORMAL_INIT_08_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_08_BIT_00_C, 1  => CPIX_NORMAL_INIT_08_BIT_01_C, 2  => CPIX_NORMAL_INIT_08_BIT_02_C, 3  => CPIX_NORMAL_INIT_08_BIT_03_C, 4  => CPIX_NORMAL_INIT_08_BIT_04_C, 5  => CPIX_NORMAL_INIT_08_BIT_05_C, 6  => CPIX_NORMAL_INIT_08_BIT_06_C, 7  => CPIX_NORMAL_INIT_08_BIT_07_C, 8  => CPIX_NORMAL_INIT_08_BIT_08_C, 9  => CPIX_NORMAL_INIT_08_BIT_09_C, 10 => CPIX_NORMAL_INIT_08_BIT_10_C, 11 => CPIX_NORMAL_INIT_08_BIT_11_C, 12 => CPIX_NORMAL_INIT_08_BIT_12_C, 13 => CPIX_NORMAL_INIT_08_BIT_13_C, 14 => CPIX_NORMAL_INIT_08_BIT_14_C);
   constant CPIX_NORMAL_INIT_09_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_09_BIT_00_C, 1  => CPIX_NORMAL_INIT_09_BIT_01_C, 2  => CPIX_NORMAL_INIT_09_BIT_02_C, 3  => CPIX_NORMAL_INIT_09_BIT_03_C, 4  => CPIX_NORMAL_INIT_09_BIT_04_C, 5  => CPIX_NORMAL_INIT_09_BIT_05_C, 6  => CPIX_NORMAL_INIT_09_BIT_06_C, 7  => CPIX_NORMAL_INIT_09_BIT_07_C, 8  => CPIX_NORMAL_INIT_09_BIT_08_C, 9  => CPIX_NORMAL_INIT_09_BIT_09_C, 10 => CPIX_NORMAL_INIT_09_BIT_10_C, 11 => CPIX_NORMAL_INIT_09_BIT_11_C, 12 => CPIX_NORMAL_INIT_09_BIT_12_C, 13 => CPIX_NORMAL_INIT_09_BIT_13_C, 14 => CPIX_NORMAL_INIT_09_BIT_14_C);
   constant CPIX_NORMAL_INIT_0A_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_0A_BIT_00_C, 1  => CPIX_NORMAL_INIT_0A_BIT_01_C, 2  => CPIX_NORMAL_INIT_0A_BIT_02_C, 3  => CPIX_NORMAL_INIT_0A_BIT_03_C, 4  => CPIX_NORMAL_INIT_0A_BIT_04_C, 5  => CPIX_NORMAL_INIT_0A_BIT_05_C, 6  => CPIX_NORMAL_INIT_0A_BIT_06_C, 7  => CPIX_NORMAL_INIT_0A_BIT_07_C, 8  => CPIX_NORMAL_INIT_0A_BIT_08_C, 9  => CPIX_NORMAL_INIT_0A_BIT_09_C, 10 => CPIX_NORMAL_INIT_0A_BIT_10_C, 11 => CPIX_NORMAL_INIT_0A_BIT_11_C, 12 => CPIX_NORMAL_INIT_0A_BIT_12_C, 13 => CPIX_NORMAL_INIT_0A_BIT_13_C, 14 => CPIX_NORMAL_INIT_0A_BIT_14_C);
   constant CPIX_NORMAL_INIT_0B_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_0B_BIT_00_C, 1  => CPIX_NORMAL_INIT_0B_BIT_01_C, 2  => CPIX_NORMAL_INIT_0B_BIT_02_C, 3  => CPIX_NORMAL_INIT_0B_BIT_03_C, 4  => CPIX_NORMAL_INIT_0B_BIT_04_C, 5  => CPIX_NORMAL_INIT_0B_BIT_05_C, 6  => CPIX_NORMAL_INIT_0B_BIT_06_C, 7  => CPIX_NORMAL_INIT_0B_BIT_07_C, 8  => CPIX_NORMAL_INIT_0B_BIT_08_C, 9  => CPIX_NORMAL_INIT_0B_BIT_09_C, 10 => CPIX_NORMAL_INIT_0B_BIT_10_C, 11 => CPIX_NORMAL_INIT_0B_BIT_11_C, 12 => CPIX_NORMAL_INIT_0B_BIT_12_C, 13 => CPIX_NORMAL_INIT_0B_BIT_13_C, 14 => CPIX_NORMAL_INIT_0B_BIT_14_C);
   constant CPIX_NORMAL_INIT_0C_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_0C_BIT_00_C, 1  => CPIX_NORMAL_INIT_0C_BIT_01_C, 2  => CPIX_NORMAL_INIT_0C_BIT_02_C, 3  => CPIX_NORMAL_INIT_0C_BIT_03_C, 4  => CPIX_NORMAL_INIT_0C_BIT_04_C, 5  => CPIX_NORMAL_INIT_0C_BIT_05_C, 6  => CPIX_NORMAL_INIT_0C_BIT_06_C, 7  => CPIX_NORMAL_INIT_0C_BIT_07_C, 8  => CPIX_NORMAL_INIT_0C_BIT_08_C, 9  => CPIX_NORMAL_INIT_0C_BIT_09_C, 10 => CPIX_NORMAL_INIT_0C_BIT_10_C, 11 => CPIX_NORMAL_INIT_0C_BIT_11_C, 12 => CPIX_NORMAL_INIT_0C_BIT_12_C, 13 => CPIX_NORMAL_INIT_0C_BIT_13_C, 14 => CPIX_NORMAL_INIT_0C_BIT_14_C);
   constant CPIX_NORMAL_INIT_0D_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_0D_BIT_00_C, 1  => CPIX_NORMAL_INIT_0D_BIT_01_C, 2  => CPIX_NORMAL_INIT_0D_BIT_02_C, 3  => CPIX_NORMAL_INIT_0D_BIT_03_C, 4  => CPIX_NORMAL_INIT_0D_BIT_04_C, 5  => CPIX_NORMAL_INIT_0D_BIT_05_C, 6  => CPIX_NORMAL_INIT_0D_BIT_06_C, 7  => CPIX_NORMAL_INIT_0D_BIT_07_C, 8  => CPIX_NORMAL_INIT_0D_BIT_08_C, 9  => CPIX_NORMAL_INIT_0D_BIT_09_C, 10 => CPIX_NORMAL_INIT_0D_BIT_10_C, 11 => CPIX_NORMAL_INIT_0D_BIT_11_C, 12 => CPIX_NORMAL_INIT_0D_BIT_12_C, 13 => CPIX_NORMAL_INIT_0D_BIT_13_C, 14 => CPIX_NORMAL_INIT_0D_BIT_14_C);
   constant CPIX_NORMAL_INIT_0E_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_0E_BIT_00_C, 1  => CPIX_NORMAL_INIT_0E_BIT_01_C, 2  => CPIX_NORMAL_INIT_0E_BIT_02_C, 3  => CPIX_NORMAL_INIT_0E_BIT_03_C, 4  => CPIX_NORMAL_INIT_0E_BIT_04_C, 5  => CPIX_NORMAL_INIT_0E_BIT_05_C, 6  => CPIX_NORMAL_INIT_0E_BIT_06_C, 7  => CPIX_NORMAL_INIT_0E_BIT_07_C, 8  => CPIX_NORMAL_INIT_0E_BIT_08_C, 9  => CPIX_NORMAL_INIT_0E_BIT_09_C, 10 => CPIX_NORMAL_INIT_0E_BIT_10_C, 11 => CPIX_NORMAL_INIT_0E_BIT_11_C, 12 => CPIX_NORMAL_INIT_0E_BIT_12_C, 13 => CPIX_NORMAL_INIT_0E_BIT_13_C, 14 => CPIX_NORMAL_INIT_0E_BIT_14_C);
   constant CPIX_NORMAL_INIT_0F_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_0F_BIT_00_C, 1  => CPIX_NORMAL_INIT_0F_BIT_01_C, 2  => CPIX_NORMAL_INIT_0F_BIT_02_C, 3  => CPIX_NORMAL_INIT_0F_BIT_03_C, 4  => CPIX_NORMAL_INIT_0F_BIT_04_C, 5  => CPIX_NORMAL_INIT_0F_BIT_05_C, 6  => CPIX_NORMAL_INIT_0F_BIT_06_C, 7  => CPIX_NORMAL_INIT_0F_BIT_07_C, 8  => CPIX_NORMAL_INIT_0F_BIT_08_C, 9  => CPIX_NORMAL_INIT_0F_BIT_09_C, 10 => CPIX_NORMAL_INIT_0F_BIT_10_C, 11 => CPIX_NORMAL_INIT_0F_BIT_11_C, 12 => CPIX_NORMAL_INIT_0F_BIT_12_C, 13 => CPIX_NORMAL_INIT_0F_BIT_13_C, 14 => CPIX_NORMAL_INIT_0F_BIT_14_C);
   constant CPIX_NORMAL_INIT_10_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_10_BIT_00_C, 1  => CPIX_NORMAL_INIT_10_BIT_01_C, 2  => CPIX_NORMAL_INIT_10_BIT_02_C, 3  => CPIX_NORMAL_INIT_10_BIT_03_C, 4  => CPIX_NORMAL_INIT_10_BIT_04_C, 5  => CPIX_NORMAL_INIT_10_BIT_05_C, 6  => CPIX_NORMAL_INIT_10_BIT_06_C, 7  => CPIX_NORMAL_INIT_10_BIT_07_C, 8  => CPIX_NORMAL_INIT_10_BIT_08_C, 9  => CPIX_NORMAL_INIT_10_BIT_09_C, 10 => CPIX_NORMAL_INIT_10_BIT_10_C, 11 => CPIX_NORMAL_INIT_10_BIT_11_C, 12 => CPIX_NORMAL_INIT_10_BIT_12_C, 13 => CPIX_NORMAL_INIT_10_BIT_13_C, 14 => CPIX_NORMAL_INIT_10_BIT_14_C);
   constant CPIX_NORMAL_INIT_11_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_11_BIT_00_C, 1  => CPIX_NORMAL_INIT_11_BIT_01_C, 2  => CPIX_NORMAL_INIT_11_BIT_02_C, 3  => CPIX_NORMAL_INIT_11_BIT_03_C, 4  => CPIX_NORMAL_INIT_11_BIT_04_C, 5  => CPIX_NORMAL_INIT_11_BIT_05_C, 6  => CPIX_NORMAL_INIT_11_BIT_06_C, 7  => CPIX_NORMAL_INIT_11_BIT_07_C, 8  => CPIX_NORMAL_INIT_11_BIT_08_C, 9  => CPIX_NORMAL_INIT_11_BIT_09_C, 10 => CPIX_NORMAL_INIT_11_BIT_10_C, 11 => CPIX_NORMAL_INIT_11_BIT_11_C, 12 => CPIX_NORMAL_INIT_11_BIT_12_C, 13 => CPIX_NORMAL_INIT_11_BIT_13_C, 14 => CPIX_NORMAL_INIT_11_BIT_14_C);
   constant CPIX_NORMAL_INIT_12_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_12_BIT_00_C, 1  => CPIX_NORMAL_INIT_12_BIT_01_C, 2  => CPIX_NORMAL_INIT_12_BIT_02_C, 3  => CPIX_NORMAL_INIT_12_BIT_03_C, 4  => CPIX_NORMAL_INIT_12_BIT_04_C, 5  => CPIX_NORMAL_INIT_12_BIT_05_C, 6  => CPIX_NORMAL_INIT_12_BIT_06_C, 7  => CPIX_NORMAL_INIT_12_BIT_07_C, 8  => CPIX_NORMAL_INIT_12_BIT_08_C, 9  => CPIX_NORMAL_INIT_12_BIT_09_C, 10 => CPIX_NORMAL_INIT_12_BIT_10_C, 11 => CPIX_NORMAL_INIT_12_BIT_11_C, 12 => CPIX_NORMAL_INIT_12_BIT_12_C, 13 => CPIX_NORMAL_INIT_12_BIT_13_C, 14 => CPIX_NORMAL_INIT_12_BIT_14_C);
   constant CPIX_NORMAL_INIT_13_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_13_BIT_00_C, 1  => CPIX_NORMAL_INIT_13_BIT_01_C, 2  => CPIX_NORMAL_INIT_13_BIT_02_C, 3  => CPIX_NORMAL_INIT_13_BIT_03_C, 4  => CPIX_NORMAL_INIT_13_BIT_04_C, 5  => CPIX_NORMAL_INIT_13_BIT_05_C, 6  => CPIX_NORMAL_INIT_13_BIT_06_C, 7  => CPIX_NORMAL_INIT_13_BIT_07_C, 8  => CPIX_NORMAL_INIT_13_BIT_08_C, 9  => CPIX_NORMAL_INIT_13_BIT_09_C, 10 => CPIX_NORMAL_INIT_13_BIT_10_C, 11 => CPIX_NORMAL_INIT_13_BIT_11_C, 12 => CPIX_NORMAL_INIT_13_BIT_12_C, 13 => CPIX_NORMAL_INIT_13_BIT_13_C, 14 => CPIX_NORMAL_INIT_13_BIT_14_C);
   constant CPIX_NORMAL_INIT_14_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_14_BIT_00_C, 1  => CPIX_NORMAL_INIT_14_BIT_01_C, 2  => CPIX_NORMAL_INIT_14_BIT_02_C, 3  => CPIX_NORMAL_INIT_14_BIT_03_C, 4  => CPIX_NORMAL_INIT_14_BIT_04_C, 5  => CPIX_NORMAL_INIT_14_BIT_05_C, 6  => CPIX_NORMAL_INIT_14_BIT_06_C, 7  => CPIX_NORMAL_INIT_14_BIT_07_C, 8  => CPIX_NORMAL_INIT_14_BIT_08_C, 9  => CPIX_NORMAL_INIT_14_BIT_09_C, 10 => CPIX_NORMAL_INIT_14_BIT_10_C, 11 => CPIX_NORMAL_INIT_14_BIT_11_C, 12 => CPIX_NORMAL_INIT_14_BIT_12_C, 13 => CPIX_NORMAL_INIT_14_BIT_13_C, 14 => CPIX_NORMAL_INIT_14_BIT_14_C);
   constant CPIX_NORMAL_INIT_15_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_15_BIT_00_C, 1  => CPIX_NORMAL_INIT_15_BIT_01_C, 2  => CPIX_NORMAL_INIT_15_BIT_02_C, 3  => CPIX_NORMAL_INIT_15_BIT_03_C, 4  => CPIX_NORMAL_INIT_15_BIT_04_C, 5  => CPIX_NORMAL_INIT_15_BIT_05_C, 6  => CPIX_NORMAL_INIT_15_BIT_06_C, 7  => CPIX_NORMAL_INIT_15_BIT_07_C, 8  => CPIX_NORMAL_INIT_15_BIT_08_C, 9  => CPIX_NORMAL_INIT_15_BIT_09_C, 10 => CPIX_NORMAL_INIT_15_BIT_10_C, 11 => CPIX_NORMAL_INIT_15_BIT_11_C, 12 => CPIX_NORMAL_INIT_15_BIT_12_C, 13 => CPIX_NORMAL_INIT_15_BIT_13_C, 14 => CPIX_NORMAL_INIT_15_BIT_14_C);
   constant CPIX_NORMAL_INIT_16_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_16_BIT_00_C, 1  => CPIX_NORMAL_INIT_16_BIT_01_C, 2  => CPIX_NORMAL_INIT_16_BIT_02_C, 3  => CPIX_NORMAL_INIT_16_BIT_03_C, 4  => CPIX_NORMAL_INIT_16_BIT_04_C, 5  => CPIX_NORMAL_INIT_16_BIT_05_C, 6  => CPIX_NORMAL_INIT_16_BIT_06_C, 7  => CPIX_NORMAL_INIT_16_BIT_07_C, 8  => CPIX_NORMAL_INIT_16_BIT_08_C, 9  => CPIX_NORMAL_INIT_16_BIT_09_C, 10 => CPIX_NORMAL_INIT_16_BIT_10_C, 11 => CPIX_NORMAL_INIT_16_BIT_11_C, 12 => CPIX_NORMAL_INIT_16_BIT_12_C, 13 => CPIX_NORMAL_INIT_16_BIT_13_C, 14 => CPIX_NORMAL_INIT_16_BIT_14_C);
   constant CPIX_NORMAL_INIT_17_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_17_BIT_00_C, 1  => CPIX_NORMAL_INIT_17_BIT_01_C, 2  => CPIX_NORMAL_INIT_17_BIT_02_C, 3  => CPIX_NORMAL_INIT_17_BIT_03_C, 4  => CPIX_NORMAL_INIT_17_BIT_04_C, 5  => CPIX_NORMAL_INIT_17_BIT_05_C, 6  => CPIX_NORMAL_INIT_17_BIT_06_C, 7  => CPIX_NORMAL_INIT_17_BIT_07_C, 8  => CPIX_NORMAL_INIT_17_BIT_08_C, 9  => CPIX_NORMAL_INIT_17_BIT_09_C, 10 => CPIX_NORMAL_INIT_17_BIT_10_C, 11 => CPIX_NORMAL_INIT_17_BIT_11_C, 12 => CPIX_NORMAL_INIT_17_BIT_12_C, 13 => CPIX_NORMAL_INIT_17_BIT_13_C, 14 => CPIX_NORMAL_INIT_17_BIT_14_C);
   constant CPIX_NORMAL_INIT_18_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_18_BIT_00_C, 1  => CPIX_NORMAL_INIT_18_BIT_01_C, 2  => CPIX_NORMAL_INIT_18_BIT_02_C, 3  => CPIX_NORMAL_INIT_18_BIT_03_C, 4  => CPIX_NORMAL_INIT_18_BIT_04_C, 5  => CPIX_NORMAL_INIT_18_BIT_05_C, 6  => CPIX_NORMAL_INIT_18_BIT_06_C, 7  => CPIX_NORMAL_INIT_18_BIT_07_C, 8  => CPIX_NORMAL_INIT_18_BIT_08_C, 9  => CPIX_NORMAL_INIT_18_BIT_09_C, 10 => CPIX_NORMAL_INIT_18_BIT_10_C, 11 => CPIX_NORMAL_INIT_18_BIT_11_C, 12 => CPIX_NORMAL_INIT_18_BIT_12_C, 13 => CPIX_NORMAL_INIT_18_BIT_13_C, 14 => CPIX_NORMAL_INIT_18_BIT_14_C);
   constant CPIX_NORMAL_INIT_19_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_19_BIT_00_C, 1  => CPIX_NORMAL_INIT_19_BIT_01_C, 2  => CPIX_NORMAL_INIT_19_BIT_02_C, 3  => CPIX_NORMAL_INIT_19_BIT_03_C, 4  => CPIX_NORMAL_INIT_19_BIT_04_C, 5  => CPIX_NORMAL_INIT_19_BIT_05_C, 6  => CPIX_NORMAL_INIT_19_BIT_06_C, 7  => CPIX_NORMAL_INIT_19_BIT_07_C, 8  => CPIX_NORMAL_INIT_19_BIT_08_C, 9  => CPIX_NORMAL_INIT_19_BIT_09_C, 10 => CPIX_NORMAL_INIT_19_BIT_10_C, 11 => CPIX_NORMAL_INIT_19_BIT_11_C, 12 => CPIX_NORMAL_INIT_19_BIT_12_C, 13 => CPIX_NORMAL_INIT_19_BIT_13_C, 14 => CPIX_NORMAL_INIT_19_BIT_14_C);
   constant CPIX_NORMAL_INIT_1A_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_1A_BIT_00_C, 1  => CPIX_NORMAL_INIT_1A_BIT_01_C, 2  => CPIX_NORMAL_INIT_1A_BIT_02_C, 3  => CPIX_NORMAL_INIT_1A_BIT_03_C, 4  => CPIX_NORMAL_INIT_1A_BIT_04_C, 5  => CPIX_NORMAL_INIT_1A_BIT_05_C, 6  => CPIX_NORMAL_INIT_1A_BIT_06_C, 7  => CPIX_NORMAL_INIT_1A_BIT_07_C, 8  => CPIX_NORMAL_INIT_1A_BIT_08_C, 9  => CPIX_NORMAL_INIT_1A_BIT_09_C, 10 => CPIX_NORMAL_INIT_1A_BIT_10_C, 11 => CPIX_NORMAL_INIT_1A_BIT_11_C, 12 => CPIX_NORMAL_INIT_1A_BIT_12_C, 13 => CPIX_NORMAL_INIT_1A_BIT_13_C, 14 => CPIX_NORMAL_INIT_1A_BIT_14_C);
   constant CPIX_NORMAL_INIT_1B_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_1B_BIT_00_C, 1  => CPIX_NORMAL_INIT_1B_BIT_01_C, 2  => CPIX_NORMAL_INIT_1B_BIT_02_C, 3  => CPIX_NORMAL_INIT_1B_BIT_03_C, 4  => CPIX_NORMAL_INIT_1B_BIT_04_C, 5  => CPIX_NORMAL_INIT_1B_BIT_05_C, 6  => CPIX_NORMAL_INIT_1B_BIT_06_C, 7  => CPIX_NORMAL_INIT_1B_BIT_07_C, 8  => CPIX_NORMAL_INIT_1B_BIT_08_C, 9  => CPIX_NORMAL_INIT_1B_BIT_09_C, 10 => CPIX_NORMAL_INIT_1B_BIT_10_C, 11 => CPIX_NORMAL_INIT_1B_BIT_11_C, 12 => CPIX_NORMAL_INIT_1B_BIT_12_C, 13 => CPIX_NORMAL_INIT_1B_BIT_13_C, 14 => CPIX_NORMAL_INIT_1B_BIT_14_C);
   constant CPIX_NORMAL_INIT_1C_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_1C_BIT_00_C, 1  => CPIX_NORMAL_INIT_1C_BIT_01_C, 2  => CPIX_NORMAL_INIT_1C_BIT_02_C, 3  => CPIX_NORMAL_INIT_1C_BIT_03_C, 4  => CPIX_NORMAL_INIT_1C_BIT_04_C, 5  => CPIX_NORMAL_INIT_1C_BIT_05_C, 6  => CPIX_NORMAL_INIT_1C_BIT_06_C, 7  => CPIX_NORMAL_INIT_1C_BIT_07_C, 8  => CPIX_NORMAL_INIT_1C_BIT_08_C, 9  => CPIX_NORMAL_INIT_1C_BIT_09_C, 10 => CPIX_NORMAL_INIT_1C_BIT_10_C, 11 => CPIX_NORMAL_INIT_1C_BIT_11_C, 12 => CPIX_NORMAL_INIT_1C_BIT_12_C, 13 => CPIX_NORMAL_INIT_1C_BIT_13_C, 14 => CPIX_NORMAL_INIT_1C_BIT_14_C);
   constant CPIX_NORMAL_INIT_1D_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_1D_BIT_00_C, 1  => CPIX_NORMAL_INIT_1D_BIT_01_C, 2  => CPIX_NORMAL_INIT_1D_BIT_02_C, 3  => CPIX_NORMAL_INIT_1D_BIT_03_C, 4  => CPIX_NORMAL_INIT_1D_BIT_04_C, 5  => CPIX_NORMAL_INIT_1D_BIT_05_C, 6  => CPIX_NORMAL_INIT_1D_BIT_06_C, 7  => CPIX_NORMAL_INIT_1D_BIT_07_C, 8  => CPIX_NORMAL_INIT_1D_BIT_08_C, 9  => CPIX_NORMAL_INIT_1D_BIT_09_C, 10 => CPIX_NORMAL_INIT_1D_BIT_10_C, 11 => CPIX_NORMAL_INIT_1D_BIT_11_C, 12 => CPIX_NORMAL_INIT_1D_BIT_12_C, 13 => CPIX_NORMAL_INIT_1D_BIT_13_C, 14 => CPIX_NORMAL_INIT_1D_BIT_14_C);
   constant CPIX_NORMAL_INIT_1E_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_1E_BIT_00_C, 1  => CPIX_NORMAL_INIT_1E_BIT_01_C, 2  => CPIX_NORMAL_INIT_1E_BIT_02_C, 3  => CPIX_NORMAL_INIT_1E_BIT_03_C, 4  => CPIX_NORMAL_INIT_1E_BIT_04_C, 5  => CPIX_NORMAL_INIT_1E_BIT_05_C, 6  => CPIX_NORMAL_INIT_1E_BIT_06_C, 7  => CPIX_NORMAL_INIT_1E_BIT_07_C, 8  => CPIX_NORMAL_INIT_1E_BIT_08_C, 9  => CPIX_NORMAL_INIT_1E_BIT_09_C, 10 => CPIX_NORMAL_INIT_1E_BIT_10_C, 11 => CPIX_NORMAL_INIT_1E_BIT_11_C, 12 => CPIX_NORMAL_INIT_1E_BIT_12_C, 13 => CPIX_NORMAL_INIT_1E_BIT_13_C, 14 => CPIX_NORMAL_INIT_1E_BIT_14_C);
   constant CPIX_NORMAL_INIT_1F_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_1F_BIT_00_C, 1  => CPIX_NORMAL_INIT_1F_BIT_01_C, 2  => CPIX_NORMAL_INIT_1F_BIT_02_C, 3  => CPIX_NORMAL_INIT_1F_BIT_03_C, 4  => CPIX_NORMAL_INIT_1F_BIT_04_C, 5  => CPIX_NORMAL_INIT_1F_BIT_05_C, 6  => CPIX_NORMAL_INIT_1F_BIT_06_C, 7  => CPIX_NORMAL_INIT_1F_BIT_07_C, 8  => CPIX_NORMAL_INIT_1F_BIT_08_C, 9  => CPIX_NORMAL_INIT_1F_BIT_09_C, 10 => CPIX_NORMAL_INIT_1F_BIT_10_C, 11 => CPIX_NORMAL_INIT_1F_BIT_11_C, 12 => CPIX_NORMAL_INIT_1F_BIT_12_C, 13 => CPIX_NORMAL_INIT_1F_BIT_13_C, 14 => CPIX_NORMAL_INIT_1F_BIT_14_C);
   constant CPIX_NORMAL_INIT_20_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_20_BIT_00_C, 1  => CPIX_NORMAL_INIT_20_BIT_01_C, 2  => CPIX_NORMAL_INIT_20_BIT_02_C, 3  => CPIX_NORMAL_INIT_20_BIT_03_C, 4  => CPIX_NORMAL_INIT_20_BIT_04_C, 5  => CPIX_NORMAL_INIT_20_BIT_05_C, 6  => CPIX_NORMAL_INIT_20_BIT_06_C, 7  => CPIX_NORMAL_INIT_20_BIT_07_C, 8  => CPIX_NORMAL_INIT_20_BIT_08_C, 9  => CPIX_NORMAL_INIT_20_BIT_09_C, 10 => CPIX_NORMAL_INIT_20_BIT_10_C, 11 => CPIX_NORMAL_INIT_20_BIT_11_C, 12 => CPIX_NORMAL_INIT_20_BIT_12_C, 13 => CPIX_NORMAL_INIT_20_BIT_13_C, 14 => CPIX_NORMAL_INIT_20_BIT_14_C);
   constant CPIX_NORMAL_INIT_21_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_21_BIT_00_C, 1  => CPIX_NORMAL_INIT_21_BIT_01_C, 2  => CPIX_NORMAL_INIT_21_BIT_02_C, 3  => CPIX_NORMAL_INIT_21_BIT_03_C, 4  => CPIX_NORMAL_INIT_21_BIT_04_C, 5  => CPIX_NORMAL_INIT_21_BIT_05_C, 6  => CPIX_NORMAL_INIT_21_BIT_06_C, 7  => CPIX_NORMAL_INIT_21_BIT_07_C, 8  => CPIX_NORMAL_INIT_21_BIT_08_C, 9  => CPIX_NORMAL_INIT_21_BIT_09_C, 10 => CPIX_NORMAL_INIT_21_BIT_10_C, 11 => CPIX_NORMAL_INIT_21_BIT_11_C, 12 => CPIX_NORMAL_INIT_21_BIT_12_C, 13 => CPIX_NORMAL_INIT_21_BIT_13_C, 14 => CPIX_NORMAL_INIT_21_BIT_14_C);
   constant CPIX_NORMAL_INIT_22_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_22_BIT_00_C, 1  => CPIX_NORMAL_INIT_22_BIT_01_C, 2  => CPIX_NORMAL_INIT_22_BIT_02_C, 3  => CPIX_NORMAL_INIT_22_BIT_03_C, 4  => CPIX_NORMAL_INIT_22_BIT_04_C, 5  => CPIX_NORMAL_INIT_22_BIT_05_C, 6  => CPIX_NORMAL_INIT_22_BIT_06_C, 7  => CPIX_NORMAL_INIT_22_BIT_07_C, 8  => CPIX_NORMAL_INIT_22_BIT_08_C, 9  => CPIX_NORMAL_INIT_22_BIT_09_C, 10 => CPIX_NORMAL_INIT_22_BIT_10_C, 11 => CPIX_NORMAL_INIT_22_BIT_11_C, 12 => CPIX_NORMAL_INIT_22_BIT_12_C, 13 => CPIX_NORMAL_INIT_22_BIT_13_C, 14 => CPIX_NORMAL_INIT_22_BIT_14_C);
   constant CPIX_NORMAL_INIT_23_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_23_BIT_00_C, 1  => CPIX_NORMAL_INIT_23_BIT_01_C, 2  => CPIX_NORMAL_INIT_23_BIT_02_C, 3  => CPIX_NORMAL_INIT_23_BIT_03_C, 4  => CPIX_NORMAL_INIT_23_BIT_04_C, 5  => CPIX_NORMAL_INIT_23_BIT_05_C, 6  => CPIX_NORMAL_INIT_23_BIT_06_C, 7  => CPIX_NORMAL_INIT_23_BIT_07_C, 8  => CPIX_NORMAL_INIT_23_BIT_08_C, 9  => CPIX_NORMAL_INIT_23_BIT_09_C, 10 => CPIX_NORMAL_INIT_23_BIT_10_C, 11 => CPIX_NORMAL_INIT_23_BIT_11_C, 12 => CPIX_NORMAL_INIT_23_BIT_12_C, 13 => CPIX_NORMAL_INIT_23_BIT_13_C, 14 => CPIX_NORMAL_INIT_23_BIT_14_C);
   constant CPIX_NORMAL_INIT_24_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_24_BIT_00_C, 1  => CPIX_NORMAL_INIT_24_BIT_01_C, 2  => CPIX_NORMAL_INIT_24_BIT_02_C, 3  => CPIX_NORMAL_INIT_24_BIT_03_C, 4  => CPIX_NORMAL_INIT_24_BIT_04_C, 5  => CPIX_NORMAL_INIT_24_BIT_05_C, 6  => CPIX_NORMAL_INIT_24_BIT_06_C, 7  => CPIX_NORMAL_INIT_24_BIT_07_C, 8  => CPIX_NORMAL_INIT_24_BIT_08_C, 9  => CPIX_NORMAL_INIT_24_BIT_09_C, 10 => CPIX_NORMAL_INIT_24_BIT_10_C, 11 => CPIX_NORMAL_INIT_24_BIT_11_C, 12 => CPIX_NORMAL_INIT_24_BIT_12_C, 13 => CPIX_NORMAL_INIT_24_BIT_13_C, 14 => CPIX_NORMAL_INIT_24_BIT_14_C);
   constant CPIX_NORMAL_INIT_25_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_25_BIT_00_C, 1  => CPIX_NORMAL_INIT_25_BIT_01_C, 2  => CPIX_NORMAL_INIT_25_BIT_02_C, 3  => CPIX_NORMAL_INIT_25_BIT_03_C, 4  => CPIX_NORMAL_INIT_25_BIT_04_C, 5  => CPIX_NORMAL_INIT_25_BIT_05_C, 6  => CPIX_NORMAL_INIT_25_BIT_06_C, 7  => CPIX_NORMAL_INIT_25_BIT_07_C, 8  => CPIX_NORMAL_INIT_25_BIT_08_C, 9  => CPIX_NORMAL_INIT_25_BIT_09_C, 10 => CPIX_NORMAL_INIT_25_BIT_10_C, 11 => CPIX_NORMAL_INIT_25_BIT_11_C, 12 => CPIX_NORMAL_INIT_25_BIT_12_C, 13 => CPIX_NORMAL_INIT_25_BIT_13_C, 14 => CPIX_NORMAL_INIT_25_BIT_14_C);
   constant CPIX_NORMAL_INIT_26_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_26_BIT_00_C, 1  => CPIX_NORMAL_INIT_26_BIT_01_C, 2  => CPIX_NORMAL_INIT_26_BIT_02_C, 3  => CPIX_NORMAL_INIT_26_BIT_03_C, 4  => CPIX_NORMAL_INIT_26_BIT_04_C, 5  => CPIX_NORMAL_INIT_26_BIT_05_C, 6  => CPIX_NORMAL_INIT_26_BIT_06_C, 7  => CPIX_NORMAL_INIT_26_BIT_07_C, 8  => CPIX_NORMAL_INIT_26_BIT_08_C, 9  => CPIX_NORMAL_INIT_26_BIT_09_C, 10 => CPIX_NORMAL_INIT_26_BIT_10_C, 11 => CPIX_NORMAL_INIT_26_BIT_11_C, 12 => CPIX_NORMAL_INIT_26_BIT_12_C, 13 => CPIX_NORMAL_INIT_26_BIT_13_C, 14 => CPIX_NORMAL_INIT_26_BIT_14_C);
   constant CPIX_NORMAL_INIT_27_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_27_BIT_00_C, 1  => CPIX_NORMAL_INIT_27_BIT_01_C, 2  => CPIX_NORMAL_INIT_27_BIT_02_C, 3  => CPIX_NORMAL_INIT_27_BIT_03_C, 4  => CPIX_NORMAL_INIT_27_BIT_04_C, 5  => CPIX_NORMAL_INIT_27_BIT_05_C, 6  => CPIX_NORMAL_INIT_27_BIT_06_C, 7  => CPIX_NORMAL_INIT_27_BIT_07_C, 8  => CPIX_NORMAL_INIT_27_BIT_08_C, 9  => CPIX_NORMAL_INIT_27_BIT_09_C, 10 => CPIX_NORMAL_INIT_27_BIT_10_C, 11 => CPIX_NORMAL_INIT_27_BIT_11_C, 12 => CPIX_NORMAL_INIT_27_BIT_12_C, 13 => CPIX_NORMAL_INIT_27_BIT_13_C, 14 => CPIX_NORMAL_INIT_27_BIT_14_C);
   constant CPIX_NORMAL_INIT_28_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_28_BIT_00_C, 1  => CPIX_NORMAL_INIT_28_BIT_01_C, 2  => CPIX_NORMAL_INIT_28_BIT_02_C, 3  => CPIX_NORMAL_INIT_28_BIT_03_C, 4  => CPIX_NORMAL_INIT_28_BIT_04_C, 5  => CPIX_NORMAL_INIT_28_BIT_05_C, 6  => CPIX_NORMAL_INIT_28_BIT_06_C, 7  => CPIX_NORMAL_INIT_28_BIT_07_C, 8  => CPIX_NORMAL_INIT_28_BIT_08_C, 9  => CPIX_NORMAL_INIT_28_BIT_09_C, 10 => CPIX_NORMAL_INIT_28_BIT_10_C, 11 => CPIX_NORMAL_INIT_28_BIT_11_C, 12 => CPIX_NORMAL_INIT_28_BIT_12_C, 13 => CPIX_NORMAL_INIT_28_BIT_13_C, 14 => CPIX_NORMAL_INIT_28_BIT_14_C);
   constant CPIX_NORMAL_INIT_29_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_29_BIT_00_C, 1  => CPIX_NORMAL_INIT_29_BIT_01_C, 2  => CPIX_NORMAL_INIT_29_BIT_02_C, 3  => CPIX_NORMAL_INIT_29_BIT_03_C, 4  => CPIX_NORMAL_INIT_29_BIT_04_C, 5  => CPIX_NORMAL_INIT_29_BIT_05_C, 6  => CPIX_NORMAL_INIT_29_BIT_06_C, 7  => CPIX_NORMAL_INIT_29_BIT_07_C, 8  => CPIX_NORMAL_INIT_29_BIT_08_C, 9  => CPIX_NORMAL_INIT_29_BIT_09_C, 10 => CPIX_NORMAL_INIT_29_BIT_10_C, 11 => CPIX_NORMAL_INIT_29_BIT_11_C, 12 => CPIX_NORMAL_INIT_29_BIT_12_C, 13 => CPIX_NORMAL_INIT_29_BIT_13_C, 14 => CPIX_NORMAL_INIT_29_BIT_14_C);
   constant CPIX_NORMAL_INIT_2A_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_2A_BIT_00_C, 1  => CPIX_NORMAL_INIT_2A_BIT_01_C, 2  => CPIX_NORMAL_INIT_2A_BIT_02_C, 3  => CPIX_NORMAL_INIT_2A_BIT_03_C, 4  => CPIX_NORMAL_INIT_2A_BIT_04_C, 5  => CPIX_NORMAL_INIT_2A_BIT_05_C, 6  => CPIX_NORMAL_INIT_2A_BIT_06_C, 7  => CPIX_NORMAL_INIT_2A_BIT_07_C, 8  => CPIX_NORMAL_INIT_2A_BIT_08_C, 9  => CPIX_NORMAL_INIT_2A_BIT_09_C, 10 => CPIX_NORMAL_INIT_2A_BIT_10_C, 11 => CPIX_NORMAL_INIT_2A_BIT_11_C, 12 => CPIX_NORMAL_INIT_2A_BIT_12_C, 13 => CPIX_NORMAL_INIT_2A_BIT_13_C, 14 => CPIX_NORMAL_INIT_2A_BIT_14_C);
   constant CPIX_NORMAL_INIT_2B_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_2B_BIT_00_C, 1  => CPIX_NORMAL_INIT_2B_BIT_01_C, 2  => CPIX_NORMAL_INIT_2B_BIT_02_C, 3  => CPIX_NORMAL_INIT_2B_BIT_03_C, 4  => CPIX_NORMAL_INIT_2B_BIT_04_C, 5  => CPIX_NORMAL_INIT_2B_BIT_05_C, 6  => CPIX_NORMAL_INIT_2B_BIT_06_C, 7  => CPIX_NORMAL_INIT_2B_BIT_07_C, 8  => CPIX_NORMAL_INIT_2B_BIT_08_C, 9  => CPIX_NORMAL_INIT_2B_BIT_09_C, 10 => CPIX_NORMAL_INIT_2B_BIT_10_C, 11 => CPIX_NORMAL_INIT_2B_BIT_11_C, 12 => CPIX_NORMAL_INIT_2B_BIT_12_C, 13 => CPIX_NORMAL_INIT_2B_BIT_13_C, 14 => CPIX_NORMAL_INIT_2B_BIT_14_C);
   constant CPIX_NORMAL_INIT_2C_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_2C_BIT_00_C, 1  => CPIX_NORMAL_INIT_2C_BIT_01_C, 2  => CPIX_NORMAL_INIT_2C_BIT_02_C, 3  => CPIX_NORMAL_INIT_2C_BIT_03_C, 4  => CPIX_NORMAL_INIT_2C_BIT_04_C, 5  => CPIX_NORMAL_INIT_2C_BIT_05_C, 6  => CPIX_NORMAL_INIT_2C_BIT_06_C, 7  => CPIX_NORMAL_INIT_2C_BIT_07_C, 8  => CPIX_NORMAL_INIT_2C_BIT_08_C, 9  => CPIX_NORMAL_INIT_2C_BIT_09_C, 10 => CPIX_NORMAL_INIT_2C_BIT_10_C, 11 => CPIX_NORMAL_INIT_2C_BIT_11_C, 12 => CPIX_NORMAL_INIT_2C_BIT_12_C, 13 => CPIX_NORMAL_INIT_2C_BIT_13_C, 14 => CPIX_NORMAL_INIT_2C_BIT_14_C);
   constant CPIX_NORMAL_INIT_2D_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_2D_BIT_00_C, 1  => CPIX_NORMAL_INIT_2D_BIT_01_C, 2  => CPIX_NORMAL_INIT_2D_BIT_02_C, 3  => CPIX_NORMAL_INIT_2D_BIT_03_C, 4  => CPIX_NORMAL_INIT_2D_BIT_04_C, 5  => CPIX_NORMAL_INIT_2D_BIT_05_C, 6  => CPIX_NORMAL_INIT_2D_BIT_06_C, 7  => CPIX_NORMAL_INIT_2D_BIT_07_C, 8  => CPIX_NORMAL_INIT_2D_BIT_08_C, 9  => CPIX_NORMAL_INIT_2D_BIT_09_C, 10 => CPIX_NORMAL_INIT_2D_BIT_10_C, 11 => CPIX_NORMAL_INIT_2D_BIT_11_C, 12 => CPIX_NORMAL_INIT_2D_BIT_12_C, 13 => CPIX_NORMAL_INIT_2D_BIT_13_C, 14 => CPIX_NORMAL_INIT_2D_BIT_14_C);
   constant CPIX_NORMAL_INIT_2E_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_2E_BIT_00_C, 1  => CPIX_NORMAL_INIT_2E_BIT_01_C, 2  => CPIX_NORMAL_INIT_2E_BIT_02_C, 3  => CPIX_NORMAL_INIT_2E_BIT_03_C, 4  => CPIX_NORMAL_INIT_2E_BIT_04_C, 5  => CPIX_NORMAL_INIT_2E_BIT_05_C, 6  => CPIX_NORMAL_INIT_2E_BIT_06_C, 7  => CPIX_NORMAL_INIT_2E_BIT_07_C, 8  => CPIX_NORMAL_INIT_2E_BIT_08_C, 9  => CPIX_NORMAL_INIT_2E_BIT_09_C, 10 => CPIX_NORMAL_INIT_2E_BIT_10_C, 11 => CPIX_NORMAL_INIT_2E_BIT_11_C, 12 => CPIX_NORMAL_INIT_2E_BIT_12_C, 13 => CPIX_NORMAL_INIT_2E_BIT_13_C, 14 => CPIX_NORMAL_INIT_2E_BIT_14_C);
   constant CPIX_NORMAL_INIT_2F_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_2F_BIT_00_C, 1  => CPIX_NORMAL_INIT_2F_BIT_01_C, 2  => CPIX_NORMAL_INIT_2F_BIT_02_C, 3  => CPIX_NORMAL_INIT_2F_BIT_03_C, 4  => CPIX_NORMAL_INIT_2F_BIT_04_C, 5  => CPIX_NORMAL_INIT_2F_BIT_05_C, 6  => CPIX_NORMAL_INIT_2F_BIT_06_C, 7  => CPIX_NORMAL_INIT_2F_BIT_07_C, 8  => CPIX_NORMAL_INIT_2F_BIT_08_C, 9  => CPIX_NORMAL_INIT_2F_BIT_09_C, 10 => CPIX_NORMAL_INIT_2F_BIT_10_C, 11 => CPIX_NORMAL_INIT_2F_BIT_11_C, 12 => CPIX_NORMAL_INIT_2F_BIT_12_C, 13 => CPIX_NORMAL_INIT_2F_BIT_13_C, 14 => CPIX_NORMAL_INIT_2F_BIT_14_C);
   constant CPIX_NORMAL_INIT_30_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_30_BIT_00_C, 1  => CPIX_NORMAL_INIT_30_BIT_01_C, 2  => CPIX_NORMAL_INIT_30_BIT_02_C, 3  => CPIX_NORMAL_INIT_30_BIT_03_C, 4  => CPIX_NORMAL_INIT_30_BIT_04_C, 5  => CPIX_NORMAL_INIT_30_BIT_05_C, 6  => CPIX_NORMAL_INIT_30_BIT_06_C, 7  => CPIX_NORMAL_INIT_30_BIT_07_C, 8  => CPIX_NORMAL_INIT_30_BIT_08_C, 9  => CPIX_NORMAL_INIT_30_BIT_09_C, 10 => CPIX_NORMAL_INIT_30_BIT_10_C, 11 => CPIX_NORMAL_INIT_30_BIT_11_C, 12 => CPIX_NORMAL_INIT_30_BIT_12_C, 13 => CPIX_NORMAL_INIT_30_BIT_13_C, 14 => CPIX_NORMAL_INIT_30_BIT_14_C);
   constant CPIX_NORMAL_INIT_31_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_31_BIT_00_C, 1  => CPIX_NORMAL_INIT_31_BIT_01_C, 2  => CPIX_NORMAL_INIT_31_BIT_02_C, 3  => CPIX_NORMAL_INIT_31_BIT_03_C, 4  => CPIX_NORMAL_INIT_31_BIT_04_C, 5  => CPIX_NORMAL_INIT_31_BIT_05_C, 6  => CPIX_NORMAL_INIT_31_BIT_06_C, 7  => CPIX_NORMAL_INIT_31_BIT_07_C, 8  => CPIX_NORMAL_INIT_31_BIT_08_C, 9  => CPIX_NORMAL_INIT_31_BIT_09_C, 10 => CPIX_NORMAL_INIT_31_BIT_10_C, 11 => CPIX_NORMAL_INIT_31_BIT_11_C, 12 => CPIX_NORMAL_INIT_31_BIT_12_C, 13 => CPIX_NORMAL_INIT_31_BIT_13_C, 14 => CPIX_NORMAL_INIT_31_BIT_14_C);
   constant CPIX_NORMAL_INIT_32_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_32_BIT_00_C, 1  => CPIX_NORMAL_INIT_32_BIT_01_C, 2  => CPIX_NORMAL_INIT_32_BIT_02_C, 3  => CPIX_NORMAL_INIT_32_BIT_03_C, 4  => CPIX_NORMAL_INIT_32_BIT_04_C, 5  => CPIX_NORMAL_INIT_32_BIT_05_C, 6  => CPIX_NORMAL_INIT_32_BIT_06_C, 7  => CPIX_NORMAL_INIT_32_BIT_07_C, 8  => CPIX_NORMAL_INIT_32_BIT_08_C, 9  => CPIX_NORMAL_INIT_32_BIT_09_C, 10 => CPIX_NORMAL_INIT_32_BIT_10_C, 11 => CPIX_NORMAL_INIT_32_BIT_11_C, 12 => CPIX_NORMAL_INIT_32_BIT_12_C, 13 => CPIX_NORMAL_INIT_32_BIT_13_C, 14 => CPIX_NORMAL_INIT_32_BIT_14_C);
   constant CPIX_NORMAL_INIT_33_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_33_BIT_00_C, 1  => CPIX_NORMAL_INIT_33_BIT_01_C, 2  => CPIX_NORMAL_INIT_33_BIT_02_C, 3  => CPIX_NORMAL_INIT_33_BIT_03_C, 4  => CPIX_NORMAL_INIT_33_BIT_04_C, 5  => CPIX_NORMAL_INIT_33_BIT_05_C, 6  => CPIX_NORMAL_INIT_33_BIT_06_C, 7  => CPIX_NORMAL_INIT_33_BIT_07_C, 8  => CPIX_NORMAL_INIT_33_BIT_08_C, 9  => CPIX_NORMAL_INIT_33_BIT_09_C, 10 => CPIX_NORMAL_INIT_33_BIT_10_C, 11 => CPIX_NORMAL_INIT_33_BIT_11_C, 12 => CPIX_NORMAL_INIT_33_BIT_12_C, 13 => CPIX_NORMAL_INIT_33_BIT_13_C, 14 => CPIX_NORMAL_INIT_33_BIT_14_C);
   constant CPIX_NORMAL_INIT_34_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_34_BIT_00_C, 1  => CPIX_NORMAL_INIT_34_BIT_01_C, 2  => CPIX_NORMAL_INIT_34_BIT_02_C, 3  => CPIX_NORMAL_INIT_34_BIT_03_C, 4  => CPIX_NORMAL_INIT_34_BIT_04_C, 5  => CPIX_NORMAL_INIT_34_BIT_05_C, 6  => CPIX_NORMAL_INIT_34_BIT_06_C, 7  => CPIX_NORMAL_INIT_34_BIT_07_C, 8  => CPIX_NORMAL_INIT_34_BIT_08_C, 9  => CPIX_NORMAL_INIT_34_BIT_09_C, 10 => CPIX_NORMAL_INIT_34_BIT_10_C, 11 => CPIX_NORMAL_INIT_34_BIT_11_C, 12 => CPIX_NORMAL_INIT_34_BIT_12_C, 13 => CPIX_NORMAL_INIT_34_BIT_13_C, 14 => CPIX_NORMAL_INIT_34_BIT_14_C);
   constant CPIX_NORMAL_INIT_35_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_35_BIT_00_C, 1  => CPIX_NORMAL_INIT_35_BIT_01_C, 2  => CPIX_NORMAL_INIT_35_BIT_02_C, 3  => CPIX_NORMAL_INIT_35_BIT_03_C, 4  => CPIX_NORMAL_INIT_35_BIT_04_C, 5  => CPIX_NORMAL_INIT_35_BIT_05_C, 6  => CPIX_NORMAL_INIT_35_BIT_06_C, 7  => CPIX_NORMAL_INIT_35_BIT_07_C, 8  => CPIX_NORMAL_INIT_35_BIT_08_C, 9  => CPIX_NORMAL_INIT_35_BIT_09_C, 10 => CPIX_NORMAL_INIT_35_BIT_10_C, 11 => CPIX_NORMAL_INIT_35_BIT_11_C, 12 => CPIX_NORMAL_INIT_35_BIT_12_C, 13 => CPIX_NORMAL_INIT_35_BIT_13_C, 14 => CPIX_NORMAL_INIT_35_BIT_14_C);
   constant CPIX_NORMAL_INIT_36_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_36_BIT_00_C, 1  => CPIX_NORMAL_INIT_36_BIT_01_C, 2  => CPIX_NORMAL_INIT_36_BIT_02_C, 3  => CPIX_NORMAL_INIT_36_BIT_03_C, 4  => CPIX_NORMAL_INIT_36_BIT_04_C, 5  => CPIX_NORMAL_INIT_36_BIT_05_C, 6  => CPIX_NORMAL_INIT_36_BIT_06_C, 7  => CPIX_NORMAL_INIT_36_BIT_07_C, 8  => CPIX_NORMAL_INIT_36_BIT_08_C, 9  => CPIX_NORMAL_INIT_36_BIT_09_C, 10 => CPIX_NORMAL_INIT_36_BIT_10_C, 11 => CPIX_NORMAL_INIT_36_BIT_11_C, 12 => CPIX_NORMAL_INIT_36_BIT_12_C, 13 => CPIX_NORMAL_INIT_36_BIT_13_C, 14 => CPIX_NORMAL_INIT_36_BIT_14_C);
   constant CPIX_NORMAL_INIT_37_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_37_BIT_00_C, 1  => CPIX_NORMAL_INIT_37_BIT_01_C, 2  => CPIX_NORMAL_INIT_37_BIT_02_C, 3  => CPIX_NORMAL_INIT_37_BIT_03_C, 4  => CPIX_NORMAL_INIT_37_BIT_04_C, 5  => CPIX_NORMAL_INIT_37_BIT_05_C, 6  => CPIX_NORMAL_INIT_37_BIT_06_C, 7  => CPIX_NORMAL_INIT_37_BIT_07_C, 8  => CPIX_NORMAL_INIT_37_BIT_08_C, 9  => CPIX_NORMAL_INIT_37_BIT_09_C, 10 => CPIX_NORMAL_INIT_37_BIT_10_C, 11 => CPIX_NORMAL_INIT_37_BIT_11_C, 12 => CPIX_NORMAL_INIT_37_BIT_12_C, 13 => CPIX_NORMAL_INIT_37_BIT_13_C, 14 => CPIX_NORMAL_INIT_37_BIT_14_C);
   constant CPIX_NORMAL_INIT_38_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_38_BIT_00_C, 1  => CPIX_NORMAL_INIT_38_BIT_01_C, 2  => CPIX_NORMAL_INIT_38_BIT_02_C, 3  => CPIX_NORMAL_INIT_38_BIT_03_C, 4  => CPIX_NORMAL_INIT_38_BIT_04_C, 5  => CPIX_NORMAL_INIT_38_BIT_05_C, 6  => CPIX_NORMAL_INIT_38_BIT_06_C, 7  => CPIX_NORMAL_INIT_38_BIT_07_C, 8  => CPIX_NORMAL_INIT_38_BIT_08_C, 9  => CPIX_NORMAL_INIT_38_BIT_09_C, 10 => CPIX_NORMAL_INIT_38_BIT_10_C, 11 => CPIX_NORMAL_INIT_38_BIT_11_C, 12 => CPIX_NORMAL_INIT_38_BIT_12_C, 13 => CPIX_NORMAL_INIT_38_BIT_13_C, 14 => CPIX_NORMAL_INIT_38_BIT_14_C);
   constant CPIX_NORMAL_INIT_39_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_39_BIT_00_C, 1  => CPIX_NORMAL_INIT_39_BIT_01_C, 2  => CPIX_NORMAL_INIT_39_BIT_02_C, 3  => CPIX_NORMAL_INIT_39_BIT_03_C, 4  => CPIX_NORMAL_INIT_39_BIT_04_C, 5  => CPIX_NORMAL_INIT_39_BIT_05_C, 6  => CPIX_NORMAL_INIT_39_BIT_06_C, 7  => CPIX_NORMAL_INIT_39_BIT_07_C, 8  => CPIX_NORMAL_INIT_39_BIT_08_C, 9  => CPIX_NORMAL_INIT_39_BIT_09_C, 10 => CPIX_NORMAL_INIT_39_BIT_10_C, 11 => CPIX_NORMAL_INIT_39_BIT_11_C, 12 => CPIX_NORMAL_INIT_39_BIT_12_C, 13 => CPIX_NORMAL_INIT_39_BIT_13_C, 14 => CPIX_NORMAL_INIT_39_BIT_14_C);
   constant CPIX_NORMAL_INIT_3A_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_3A_BIT_00_C, 1  => CPIX_NORMAL_INIT_3A_BIT_01_C, 2  => CPIX_NORMAL_INIT_3A_BIT_02_C, 3  => CPIX_NORMAL_INIT_3A_BIT_03_C, 4  => CPIX_NORMAL_INIT_3A_BIT_04_C, 5  => CPIX_NORMAL_INIT_3A_BIT_05_C, 6  => CPIX_NORMAL_INIT_3A_BIT_06_C, 7  => CPIX_NORMAL_INIT_3A_BIT_07_C, 8  => CPIX_NORMAL_INIT_3A_BIT_08_C, 9  => CPIX_NORMAL_INIT_3A_BIT_09_C, 10 => CPIX_NORMAL_INIT_3A_BIT_10_C, 11 => CPIX_NORMAL_INIT_3A_BIT_11_C, 12 => CPIX_NORMAL_INIT_3A_BIT_12_C, 13 => CPIX_NORMAL_INIT_3A_BIT_13_C, 14 => CPIX_NORMAL_INIT_3A_BIT_14_C);
   constant CPIX_NORMAL_INIT_3B_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_3B_BIT_00_C, 1  => CPIX_NORMAL_INIT_3B_BIT_01_C, 2  => CPIX_NORMAL_INIT_3B_BIT_02_C, 3  => CPIX_NORMAL_INIT_3B_BIT_03_C, 4  => CPIX_NORMAL_INIT_3B_BIT_04_C, 5  => CPIX_NORMAL_INIT_3B_BIT_05_C, 6  => CPIX_NORMAL_INIT_3B_BIT_06_C, 7  => CPIX_NORMAL_INIT_3B_BIT_07_C, 8  => CPIX_NORMAL_INIT_3B_BIT_08_C, 9  => CPIX_NORMAL_INIT_3B_BIT_09_C, 10 => CPIX_NORMAL_INIT_3B_BIT_10_C, 11 => CPIX_NORMAL_INIT_3B_BIT_11_C, 12 => CPIX_NORMAL_INIT_3B_BIT_12_C, 13 => CPIX_NORMAL_INIT_3B_BIT_13_C, 14 => CPIX_NORMAL_INIT_3B_BIT_14_C);
   constant CPIX_NORMAL_INIT_3C_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_3C_BIT_00_C, 1  => CPIX_NORMAL_INIT_3C_BIT_01_C, 2  => CPIX_NORMAL_INIT_3C_BIT_02_C, 3  => CPIX_NORMAL_INIT_3C_BIT_03_C, 4  => CPIX_NORMAL_INIT_3C_BIT_04_C, 5  => CPIX_NORMAL_INIT_3C_BIT_05_C, 6  => CPIX_NORMAL_INIT_3C_BIT_06_C, 7  => CPIX_NORMAL_INIT_3C_BIT_07_C, 8  => CPIX_NORMAL_INIT_3C_BIT_08_C, 9  => CPIX_NORMAL_INIT_3C_BIT_09_C, 10 => CPIX_NORMAL_INIT_3C_BIT_10_C, 11 => CPIX_NORMAL_INIT_3C_BIT_11_C, 12 => CPIX_NORMAL_INIT_3C_BIT_12_C, 13 => CPIX_NORMAL_INIT_3C_BIT_13_C, 14 => CPIX_NORMAL_INIT_3C_BIT_14_C);
   constant CPIX_NORMAL_INIT_3D_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_3D_BIT_00_C, 1  => CPIX_NORMAL_INIT_3D_BIT_01_C, 2  => CPIX_NORMAL_INIT_3D_BIT_02_C, 3  => CPIX_NORMAL_INIT_3D_BIT_03_C, 4  => CPIX_NORMAL_INIT_3D_BIT_04_C, 5  => CPIX_NORMAL_INIT_3D_BIT_05_C, 6  => CPIX_NORMAL_INIT_3D_BIT_06_C, 7  => CPIX_NORMAL_INIT_3D_BIT_07_C, 8  => CPIX_NORMAL_INIT_3D_BIT_08_C, 9  => CPIX_NORMAL_INIT_3D_BIT_09_C, 10 => CPIX_NORMAL_INIT_3D_BIT_10_C, 11 => CPIX_NORMAL_INIT_3D_BIT_11_C, 12 => CPIX_NORMAL_INIT_3D_BIT_12_C, 13 => CPIX_NORMAL_INIT_3D_BIT_13_C, 14 => CPIX_NORMAL_INIT_3D_BIT_14_C);
   constant CPIX_NORMAL_INIT_3E_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_3E_BIT_00_C, 1  => CPIX_NORMAL_INIT_3E_BIT_01_C, 2  => CPIX_NORMAL_INIT_3E_BIT_02_C, 3  => CPIX_NORMAL_INIT_3E_BIT_03_C, 4  => CPIX_NORMAL_INIT_3E_BIT_04_C, 5  => CPIX_NORMAL_INIT_3E_BIT_05_C, 6  => CPIX_NORMAL_INIT_3E_BIT_06_C, 7  => CPIX_NORMAL_INIT_3E_BIT_07_C, 8  => CPIX_NORMAL_INIT_3E_BIT_08_C, 9  => CPIX_NORMAL_INIT_3E_BIT_09_C, 10 => CPIX_NORMAL_INIT_3E_BIT_10_C, 11 => CPIX_NORMAL_INIT_3E_BIT_11_C, 12 => CPIX_NORMAL_INIT_3E_BIT_12_C, 13 => CPIX_NORMAL_INIT_3E_BIT_13_C, 14 => CPIX_NORMAL_INIT_3E_BIT_14_C);
   constant CPIX_NORMAL_INIT_3F_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_3F_BIT_00_C, 1  => CPIX_NORMAL_INIT_3F_BIT_01_C, 2  => CPIX_NORMAL_INIT_3F_BIT_02_C, 3  => CPIX_NORMAL_INIT_3F_BIT_03_C, 4  => CPIX_NORMAL_INIT_3F_BIT_04_C, 5  => CPIX_NORMAL_INIT_3F_BIT_05_C, 6  => CPIX_NORMAL_INIT_3F_BIT_06_C, 7  => CPIX_NORMAL_INIT_3F_BIT_07_C, 8  => CPIX_NORMAL_INIT_3F_BIT_08_C, 9  => CPIX_NORMAL_INIT_3F_BIT_09_C, 10 => CPIX_NORMAL_INIT_3F_BIT_10_C, 11 => CPIX_NORMAL_INIT_3F_BIT_11_C, 12 => CPIX_NORMAL_INIT_3F_BIT_12_C, 13 => CPIX_NORMAL_INIT_3F_BIT_13_C, 14 => CPIX_NORMAL_INIT_3F_BIT_14_C);
   constant CPIX_NORMAL_INIT_40_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_40_BIT_00_C, 1  => CPIX_NORMAL_INIT_40_BIT_01_C, 2  => CPIX_NORMAL_INIT_40_BIT_02_C, 3  => CPIX_NORMAL_INIT_40_BIT_03_C, 4  => CPIX_NORMAL_INIT_40_BIT_04_C, 5  => CPIX_NORMAL_INIT_40_BIT_05_C, 6  => CPIX_NORMAL_INIT_40_BIT_06_C, 7  => CPIX_NORMAL_INIT_40_BIT_07_C, 8  => CPIX_NORMAL_INIT_40_BIT_08_C, 9  => CPIX_NORMAL_INIT_40_BIT_09_C, 10 => CPIX_NORMAL_INIT_40_BIT_10_C, 11 => CPIX_NORMAL_INIT_40_BIT_11_C, 12 => CPIX_NORMAL_INIT_40_BIT_12_C, 13 => CPIX_NORMAL_INIT_40_BIT_13_C, 14 => CPIX_NORMAL_INIT_40_BIT_14_C);
   constant CPIX_NORMAL_INIT_41_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_41_BIT_00_C, 1  => CPIX_NORMAL_INIT_41_BIT_01_C, 2  => CPIX_NORMAL_INIT_41_BIT_02_C, 3  => CPIX_NORMAL_INIT_41_BIT_03_C, 4  => CPIX_NORMAL_INIT_41_BIT_04_C, 5  => CPIX_NORMAL_INIT_41_BIT_05_C, 6  => CPIX_NORMAL_INIT_41_BIT_06_C, 7  => CPIX_NORMAL_INIT_41_BIT_07_C, 8  => CPIX_NORMAL_INIT_41_BIT_08_C, 9  => CPIX_NORMAL_INIT_41_BIT_09_C, 10 => CPIX_NORMAL_INIT_41_BIT_10_C, 11 => CPIX_NORMAL_INIT_41_BIT_11_C, 12 => CPIX_NORMAL_INIT_41_BIT_12_C, 13 => CPIX_NORMAL_INIT_41_BIT_13_C, 14 => CPIX_NORMAL_INIT_41_BIT_14_C);
   constant CPIX_NORMAL_INIT_42_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_42_BIT_00_C, 1  => CPIX_NORMAL_INIT_42_BIT_01_C, 2  => CPIX_NORMAL_INIT_42_BIT_02_C, 3  => CPIX_NORMAL_INIT_42_BIT_03_C, 4  => CPIX_NORMAL_INIT_42_BIT_04_C, 5  => CPIX_NORMAL_INIT_42_BIT_05_C, 6  => CPIX_NORMAL_INIT_42_BIT_06_C, 7  => CPIX_NORMAL_INIT_42_BIT_07_C, 8  => CPIX_NORMAL_INIT_42_BIT_08_C, 9  => CPIX_NORMAL_INIT_42_BIT_09_C, 10 => CPIX_NORMAL_INIT_42_BIT_10_C, 11 => CPIX_NORMAL_INIT_42_BIT_11_C, 12 => CPIX_NORMAL_INIT_42_BIT_12_C, 13 => CPIX_NORMAL_INIT_42_BIT_13_C, 14 => CPIX_NORMAL_INIT_42_BIT_14_C);
   constant CPIX_NORMAL_INIT_43_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_43_BIT_00_C, 1  => CPIX_NORMAL_INIT_43_BIT_01_C, 2  => CPIX_NORMAL_INIT_43_BIT_02_C, 3  => CPIX_NORMAL_INIT_43_BIT_03_C, 4  => CPIX_NORMAL_INIT_43_BIT_04_C, 5  => CPIX_NORMAL_INIT_43_BIT_05_C, 6  => CPIX_NORMAL_INIT_43_BIT_06_C, 7  => CPIX_NORMAL_INIT_43_BIT_07_C, 8  => CPIX_NORMAL_INIT_43_BIT_08_C, 9  => CPIX_NORMAL_INIT_43_BIT_09_C, 10 => CPIX_NORMAL_INIT_43_BIT_10_C, 11 => CPIX_NORMAL_INIT_43_BIT_11_C, 12 => CPIX_NORMAL_INIT_43_BIT_12_C, 13 => CPIX_NORMAL_INIT_43_BIT_13_C, 14 => CPIX_NORMAL_INIT_43_BIT_14_C);
   constant CPIX_NORMAL_INIT_44_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_44_BIT_00_C, 1  => CPIX_NORMAL_INIT_44_BIT_01_C, 2  => CPIX_NORMAL_INIT_44_BIT_02_C, 3  => CPIX_NORMAL_INIT_44_BIT_03_C, 4  => CPIX_NORMAL_INIT_44_BIT_04_C, 5  => CPIX_NORMAL_INIT_44_BIT_05_C, 6  => CPIX_NORMAL_INIT_44_BIT_06_C, 7  => CPIX_NORMAL_INIT_44_BIT_07_C, 8  => CPIX_NORMAL_INIT_44_BIT_08_C, 9  => CPIX_NORMAL_INIT_44_BIT_09_C, 10 => CPIX_NORMAL_INIT_44_BIT_10_C, 11 => CPIX_NORMAL_INIT_44_BIT_11_C, 12 => CPIX_NORMAL_INIT_44_BIT_12_C, 13 => CPIX_NORMAL_INIT_44_BIT_13_C, 14 => CPIX_NORMAL_INIT_44_BIT_14_C);
   constant CPIX_NORMAL_INIT_45_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_45_BIT_00_C, 1  => CPIX_NORMAL_INIT_45_BIT_01_C, 2  => CPIX_NORMAL_INIT_45_BIT_02_C, 3  => CPIX_NORMAL_INIT_45_BIT_03_C, 4  => CPIX_NORMAL_INIT_45_BIT_04_C, 5  => CPIX_NORMAL_INIT_45_BIT_05_C, 6  => CPIX_NORMAL_INIT_45_BIT_06_C, 7  => CPIX_NORMAL_INIT_45_BIT_07_C, 8  => CPIX_NORMAL_INIT_45_BIT_08_C, 9  => CPIX_NORMAL_INIT_45_BIT_09_C, 10 => CPIX_NORMAL_INIT_45_BIT_10_C, 11 => CPIX_NORMAL_INIT_45_BIT_11_C, 12 => CPIX_NORMAL_INIT_45_BIT_12_C, 13 => CPIX_NORMAL_INIT_45_BIT_13_C, 14 => CPIX_NORMAL_INIT_45_BIT_14_C);
   constant CPIX_NORMAL_INIT_46_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_46_BIT_00_C, 1  => CPIX_NORMAL_INIT_46_BIT_01_C, 2  => CPIX_NORMAL_INIT_46_BIT_02_C, 3  => CPIX_NORMAL_INIT_46_BIT_03_C, 4  => CPIX_NORMAL_INIT_46_BIT_04_C, 5  => CPIX_NORMAL_INIT_46_BIT_05_C, 6  => CPIX_NORMAL_INIT_46_BIT_06_C, 7  => CPIX_NORMAL_INIT_46_BIT_07_C, 8  => CPIX_NORMAL_INIT_46_BIT_08_C, 9  => CPIX_NORMAL_INIT_46_BIT_09_C, 10 => CPIX_NORMAL_INIT_46_BIT_10_C, 11 => CPIX_NORMAL_INIT_46_BIT_11_C, 12 => CPIX_NORMAL_INIT_46_BIT_12_C, 13 => CPIX_NORMAL_INIT_46_BIT_13_C, 14 => CPIX_NORMAL_INIT_46_BIT_14_C);
   constant CPIX_NORMAL_INIT_47_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_47_BIT_00_C, 1  => CPIX_NORMAL_INIT_47_BIT_01_C, 2  => CPIX_NORMAL_INIT_47_BIT_02_C, 3  => CPIX_NORMAL_INIT_47_BIT_03_C, 4  => CPIX_NORMAL_INIT_47_BIT_04_C, 5  => CPIX_NORMAL_INIT_47_BIT_05_C, 6  => CPIX_NORMAL_INIT_47_BIT_06_C, 7  => CPIX_NORMAL_INIT_47_BIT_07_C, 8  => CPIX_NORMAL_INIT_47_BIT_08_C, 9  => CPIX_NORMAL_INIT_47_BIT_09_C, 10 => CPIX_NORMAL_INIT_47_BIT_10_C, 11 => CPIX_NORMAL_INIT_47_BIT_11_C, 12 => CPIX_NORMAL_INIT_47_BIT_12_C, 13 => CPIX_NORMAL_INIT_47_BIT_13_C, 14 => CPIX_NORMAL_INIT_47_BIT_14_C);
   constant CPIX_NORMAL_INIT_48_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_48_BIT_00_C, 1  => CPIX_NORMAL_INIT_48_BIT_01_C, 2  => CPIX_NORMAL_INIT_48_BIT_02_C, 3  => CPIX_NORMAL_INIT_48_BIT_03_C, 4  => CPIX_NORMAL_INIT_48_BIT_04_C, 5  => CPIX_NORMAL_INIT_48_BIT_05_C, 6  => CPIX_NORMAL_INIT_48_BIT_06_C, 7  => CPIX_NORMAL_INIT_48_BIT_07_C, 8  => CPIX_NORMAL_INIT_48_BIT_08_C, 9  => CPIX_NORMAL_INIT_48_BIT_09_C, 10 => CPIX_NORMAL_INIT_48_BIT_10_C, 11 => CPIX_NORMAL_INIT_48_BIT_11_C, 12 => CPIX_NORMAL_INIT_48_BIT_12_C, 13 => CPIX_NORMAL_INIT_48_BIT_13_C, 14 => CPIX_NORMAL_INIT_48_BIT_14_C);
   constant CPIX_NORMAL_INIT_49_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_49_BIT_00_C, 1  => CPIX_NORMAL_INIT_49_BIT_01_C, 2  => CPIX_NORMAL_INIT_49_BIT_02_C, 3  => CPIX_NORMAL_INIT_49_BIT_03_C, 4  => CPIX_NORMAL_INIT_49_BIT_04_C, 5  => CPIX_NORMAL_INIT_49_BIT_05_C, 6  => CPIX_NORMAL_INIT_49_BIT_06_C, 7  => CPIX_NORMAL_INIT_49_BIT_07_C, 8  => CPIX_NORMAL_INIT_49_BIT_08_C, 9  => CPIX_NORMAL_INIT_49_BIT_09_C, 10 => CPIX_NORMAL_INIT_49_BIT_10_C, 11 => CPIX_NORMAL_INIT_49_BIT_11_C, 12 => CPIX_NORMAL_INIT_49_BIT_12_C, 13 => CPIX_NORMAL_INIT_49_BIT_13_C, 14 => CPIX_NORMAL_INIT_49_BIT_14_C);
   constant CPIX_NORMAL_INIT_4A_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_4A_BIT_00_C, 1  => CPIX_NORMAL_INIT_4A_BIT_01_C, 2  => CPIX_NORMAL_INIT_4A_BIT_02_C, 3  => CPIX_NORMAL_INIT_4A_BIT_03_C, 4  => CPIX_NORMAL_INIT_4A_BIT_04_C, 5  => CPIX_NORMAL_INIT_4A_BIT_05_C, 6  => CPIX_NORMAL_INIT_4A_BIT_06_C, 7  => CPIX_NORMAL_INIT_4A_BIT_07_C, 8  => CPIX_NORMAL_INIT_4A_BIT_08_C, 9  => CPIX_NORMAL_INIT_4A_BIT_09_C, 10 => CPIX_NORMAL_INIT_4A_BIT_10_C, 11 => CPIX_NORMAL_INIT_4A_BIT_11_C, 12 => CPIX_NORMAL_INIT_4A_BIT_12_C, 13 => CPIX_NORMAL_INIT_4A_BIT_13_C, 14 => CPIX_NORMAL_INIT_4A_BIT_14_C);
   constant CPIX_NORMAL_INIT_4B_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_4B_BIT_00_C, 1  => CPIX_NORMAL_INIT_4B_BIT_01_C, 2  => CPIX_NORMAL_INIT_4B_BIT_02_C, 3  => CPIX_NORMAL_INIT_4B_BIT_03_C, 4  => CPIX_NORMAL_INIT_4B_BIT_04_C, 5  => CPIX_NORMAL_INIT_4B_BIT_05_C, 6  => CPIX_NORMAL_INIT_4B_BIT_06_C, 7  => CPIX_NORMAL_INIT_4B_BIT_07_C, 8  => CPIX_NORMAL_INIT_4B_BIT_08_C, 9  => CPIX_NORMAL_INIT_4B_BIT_09_C, 10 => CPIX_NORMAL_INIT_4B_BIT_10_C, 11 => CPIX_NORMAL_INIT_4B_BIT_11_C, 12 => CPIX_NORMAL_INIT_4B_BIT_12_C, 13 => CPIX_NORMAL_INIT_4B_BIT_13_C, 14 => CPIX_NORMAL_INIT_4B_BIT_14_C);
   constant CPIX_NORMAL_INIT_4C_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_4C_BIT_00_C, 1  => CPIX_NORMAL_INIT_4C_BIT_01_C, 2  => CPIX_NORMAL_INIT_4C_BIT_02_C, 3  => CPIX_NORMAL_INIT_4C_BIT_03_C, 4  => CPIX_NORMAL_INIT_4C_BIT_04_C, 5  => CPIX_NORMAL_INIT_4C_BIT_05_C, 6  => CPIX_NORMAL_INIT_4C_BIT_06_C, 7  => CPIX_NORMAL_INIT_4C_BIT_07_C, 8  => CPIX_NORMAL_INIT_4C_BIT_08_C, 9  => CPIX_NORMAL_INIT_4C_BIT_09_C, 10 => CPIX_NORMAL_INIT_4C_BIT_10_C, 11 => CPIX_NORMAL_INIT_4C_BIT_11_C, 12 => CPIX_NORMAL_INIT_4C_BIT_12_C, 13 => CPIX_NORMAL_INIT_4C_BIT_13_C, 14 => CPIX_NORMAL_INIT_4C_BIT_14_C);
   constant CPIX_NORMAL_INIT_4D_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_4D_BIT_00_C, 1  => CPIX_NORMAL_INIT_4D_BIT_01_C, 2  => CPIX_NORMAL_INIT_4D_BIT_02_C, 3  => CPIX_NORMAL_INIT_4D_BIT_03_C, 4  => CPIX_NORMAL_INIT_4D_BIT_04_C, 5  => CPIX_NORMAL_INIT_4D_BIT_05_C, 6  => CPIX_NORMAL_INIT_4D_BIT_06_C, 7  => CPIX_NORMAL_INIT_4D_BIT_07_C, 8  => CPIX_NORMAL_INIT_4D_BIT_08_C, 9  => CPIX_NORMAL_INIT_4D_BIT_09_C, 10 => CPIX_NORMAL_INIT_4D_BIT_10_C, 11 => CPIX_NORMAL_INIT_4D_BIT_11_C, 12 => CPIX_NORMAL_INIT_4D_BIT_12_C, 13 => CPIX_NORMAL_INIT_4D_BIT_13_C, 14 => CPIX_NORMAL_INIT_4D_BIT_14_C);
   constant CPIX_NORMAL_INIT_4E_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_4E_BIT_00_C, 1  => CPIX_NORMAL_INIT_4E_BIT_01_C, 2  => CPIX_NORMAL_INIT_4E_BIT_02_C, 3  => CPIX_NORMAL_INIT_4E_BIT_03_C, 4  => CPIX_NORMAL_INIT_4E_BIT_04_C, 5  => CPIX_NORMAL_INIT_4E_BIT_05_C, 6  => CPIX_NORMAL_INIT_4E_BIT_06_C, 7  => CPIX_NORMAL_INIT_4E_BIT_07_C, 8  => CPIX_NORMAL_INIT_4E_BIT_08_C, 9  => CPIX_NORMAL_INIT_4E_BIT_09_C, 10 => CPIX_NORMAL_INIT_4E_BIT_10_C, 11 => CPIX_NORMAL_INIT_4E_BIT_11_C, 12 => CPIX_NORMAL_INIT_4E_BIT_12_C, 13 => CPIX_NORMAL_INIT_4E_BIT_13_C, 14 => CPIX_NORMAL_INIT_4E_BIT_14_C);
   constant CPIX_NORMAL_INIT_4F_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_4F_BIT_00_C, 1  => CPIX_NORMAL_INIT_4F_BIT_01_C, 2  => CPIX_NORMAL_INIT_4F_BIT_02_C, 3  => CPIX_NORMAL_INIT_4F_BIT_03_C, 4  => CPIX_NORMAL_INIT_4F_BIT_04_C, 5  => CPIX_NORMAL_INIT_4F_BIT_05_C, 6  => CPIX_NORMAL_INIT_4F_BIT_06_C, 7  => CPIX_NORMAL_INIT_4F_BIT_07_C, 8  => CPIX_NORMAL_INIT_4F_BIT_08_C, 9  => CPIX_NORMAL_INIT_4F_BIT_09_C, 10 => CPIX_NORMAL_INIT_4F_BIT_10_C, 11 => CPIX_NORMAL_INIT_4F_BIT_11_C, 12 => CPIX_NORMAL_INIT_4F_BIT_12_C, 13 => CPIX_NORMAL_INIT_4F_BIT_13_C, 14 => CPIX_NORMAL_INIT_4F_BIT_14_C);
   constant CPIX_NORMAL_INIT_50_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_50_BIT_00_C, 1  => CPIX_NORMAL_INIT_50_BIT_01_C, 2  => CPIX_NORMAL_INIT_50_BIT_02_C, 3  => CPIX_NORMAL_INIT_50_BIT_03_C, 4  => CPIX_NORMAL_INIT_50_BIT_04_C, 5  => CPIX_NORMAL_INIT_50_BIT_05_C, 6  => CPIX_NORMAL_INIT_50_BIT_06_C, 7  => CPIX_NORMAL_INIT_50_BIT_07_C, 8  => CPIX_NORMAL_INIT_50_BIT_08_C, 9  => CPIX_NORMAL_INIT_50_BIT_09_C, 10 => CPIX_NORMAL_INIT_50_BIT_10_C, 11 => CPIX_NORMAL_INIT_50_BIT_11_C, 12 => CPIX_NORMAL_INIT_50_BIT_12_C, 13 => CPIX_NORMAL_INIT_50_BIT_13_C, 14 => CPIX_NORMAL_INIT_50_BIT_14_C);
   constant CPIX_NORMAL_INIT_51_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_51_BIT_00_C, 1  => CPIX_NORMAL_INIT_51_BIT_01_C, 2  => CPIX_NORMAL_INIT_51_BIT_02_C, 3  => CPIX_NORMAL_INIT_51_BIT_03_C, 4  => CPIX_NORMAL_INIT_51_BIT_04_C, 5  => CPIX_NORMAL_INIT_51_BIT_05_C, 6  => CPIX_NORMAL_INIT_51_BIT_06_C, 7  => CPIX_NORMAL_INIT_51_BIT_07_C, 8  => CPIX_NORMAL_INIT_51_BIT_08_C, 9  => CPIX_NORMAL_INIT_51_BIT_09_C, 10 => CPIX_NORMAL_INIT_51_BIT_10_C, 11 => CPIX_NORMAL_INIT_51_BIT_11_C, 12 => CPIX_NORMAL_INIT_51_BIT_12_C, 13 => CPIX_NORMAL_INIT_51_BIT_13_C, 14 => CPIX_NORMAL_INIT_51_BIT_14_C);
   constant CPIX_NORMAL_INIT_52_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_52_BIT_00_C, 1  => CPIX_NORMAL_INIT_52_BIT_01_C, 2  => CPIX_NORMAL_INIT_52_BIT_02_C, 3  => CPIX_NORMAL_INIT_52_BIT_03_C, 4  => CPIX_NORMAL_INIT_52_BIT_04_C, 5  => CPIX_NORMAL_INIT_52_BIT_05_C, 6  => CPIX_NORMAL_INIT_52_BIT_06_C, 7  => CPIX_NORMAL_INIT_52_BIT_07_C, 8  => CPIX_NORMAL_INIT_52_BIT_08_C, 9  => CPIX_NORMAL_INIT_52_BIT_09_C, 10 => CPIX_NORMAL_INIT_52_BIT_10_C, 11 => CPIX_NORMAL_INIT_52_BIT_11_C, 12 => CPIX_NORMAL_INIT_52_BIT_12_C, 13 => CPIX_NORMAL_INIT_52_BIT_13_C, 14 => CPIX_NORMAL_INIT_52_BIT_14_C);
   constant CPIX_NORMAL_INIT_53_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_53_BIT_00_C, 1  => CPIX_NORMAL_INIT_53_BIT_01_C, 2  => CPIX_NORMAL_INIT_53_BIT_02_C, 3  => CPIX_NORMAL_INIT_53_BIT_03_C, 4  => CPIX_NORMAL_INIT_53_BIT_04_C, 5  => CPIX_NORMAL_INIT_53_BIT_05_C, 6  => CPIX_NORMAL_INIT_53_BIT_06_C, 7  => CPIX_NORMAL_INIT_53_BIT_07_C, 8  => CPIX_NORMAL_INIT_53_BIT_08_C, 9  => CPIX_NORMAL_INIT_53_BIT_09_C, 10 => CPIX_NORMAL_INIT_53_BIT_10_C, 11 => CPIX_NORMAL_INIT_53_BIT_11_C, 12 => CPIX_NORMAL_INIT_53_BIT_12_C, 13 => CPIX_NORMAL_INIT_53_BIT_13_C, 14 => CPIX_NORMAL_INIT_53_BIT_14_C);
   constant CPIX_NORMAL_INIT_54_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_54_BIT_00_C, 1  => CPIX_NORMAL_INIT_54_BIT_01_C, 2  => CPIX_NORMAL_INIT_54_BIT_02_C, 3  => CPIX_NORMAL_INIT_54_BIT_03_C, 4  => CPIX_NORMAL_INIT_54_BIT_04_C, 5  => CPIX_NORMAL_INIT_54_BIT_05_C, 6  => CPIX_NORMAL_INIT_54_BIT_06_C, 7  => CPIX_NORMAL_INIT_54_BIT_07_C, 8  => CPIX_NORMAL_INIT_54_BIT_08_C, 9  => CPIX_NORMAL_INIT_54_BIT_09_C, 10 => CPIX_NORMAL_INIT_54_BIT_10_C, 11 => CPIX_NORMAL_INIT_54_BIT_11_C, 12 => CPIX_NORMAL_INIT_54_BIT_12_C, 13 => CPIX_NORMAL_INIT_54_BIT_13_C, 14 => CPIX_NORMAL_INIT_54_BIT_14_C);
   constant CPIX_NORMAL_INIT_55_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_55_BIT_00_C, 1  => CPIX_NORMAL_INIT_55_BIT_01_C, 2  => CPIX_NORMAL_INIT_55_BIT_02_C, 3  => CPIX_NORMAL_INIT_55_BIT_03_C, 4  => CPIX_NORMAL_INIT_55_BIT_04_C, 5  => CPIX_NORMAL_INIT_55_BIT_05_C, 6  => CPIX_NORMAL_INIT_55_BIT_06_C, 7  => CPIX_NORMAL_INIT_55_BIT_07_C, 8  => CPIX_NORMAL_INIT_55_BIT_08_C, 9  => CPIX_NORMAL_INIT_55_BIT_09_C, 10 => CPIX_NORMAL_INIT_55_BIT_10_C, 11 => CPIX_NORMAL_INIT_55_BIT_11_C, 12 => CPIX_NORMAL_INIT_55_BIT_12_C, 13 => CPIX_NORMAL_INIT_55_BIT_13_C, 14 => CPIX_NORMAL_INIT_55_BIT_14_C);
   constant CPIX_NORMAL_INIT_56_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_56_BIT_00_C, 1  => CPIX_NORMAL_INIT_56_BIT_01_C, 2  => CPIX_NORMAL_INIT_56_BIT_02_C, 3  => CPIX_NORMAL_INIT_56_BIT_03_C, 4  => CPIX_NORMAL_INIT_56_BIT_04_C, 5  => CPIX_NORMAL_INIT_56_BIT_05_C, 6  => CPIX_NORMAL_INIT_56_BIT_06_C, 7  => CPIX_NORMAL_INIT_56_BIT_07_C, 8  => CPIX_NORMAL_INIT_56_BIT_08_C, 9  => CPIX_NORMAL_INIT_56_BIT_09_C, 10 => CPIX_NORMAL_INIT_56_BIT_10_C, 11 => CPIX_NORMAL_INIT_56_BIT_11_C, 12 => CPIX_NORMAL_INIT_56_BIT_12_C, 13 => CPIX_NORMAL_INIT_56_BIT_13_C, 14 => CPIX_NORMAL_INIT_56_BIT_14_C);
   constant CPIX_NORMAL_INIT_57_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_57_BIT_00_C, 1  => CPIX_NORMAL_INIT_57_BIT_01_C, 2  => CPIX_NORMAL_INIT_57_BIT_02_C, 3  => CPIX_NORMAL_INIT_57_BIT_03_C, 4  => CPIX_NORMAL_INIT_57_BIT_04_C, 5  => CPIX_NORMAL_INIT_57_BIT_05_C, 6  => CPIX_NORMAL_INIT_57_BIT_06_C, 7  => CPIX_NORMAL_INIT_57_BIT_07_C, 8  => CPIX_NORMAL_INIT_57_BIT_08_C, 9  => CPIX_NORMAL_INIT_57_BIT_09_C, 10 => CPIX_NORMAL_INIT_57_BIT_10_C, 11 => CPIX_NORMAL_INIT_57_BIT_11_C, 12 => CPIX_NORMAL_INIT_57_BIT_12_C, 13 => CPIX_NORMAL_INIT_57_BIT_13_C, 14 => CPIX_NORMAL_INIT_57_BIT_14_C);
   constant CPIX_NORMAL_INIT_58_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_58_BIT_00_C, 1  => CPIX_NORMAL_INIT_58_BIT_01_C, 2  => CPIX_NORMAL_INIT_58_BIT_02_C, 3  => CPIX_NORMAL_INIT_58_BIT_03_C, 4  => CPIX_NORMAL_INIT_58_BIT_04_C, 5  => CPIX_NORMAL_INIT_58_BIT_05_C, 6  => CPIX_NORMAL_INIT_58_BIT_06_C, 7  => CPIX_NORMAL_INIT_58_BIT_07_C, 8  => CPIX_NORMAL_INIT_58_BIT_08_C, 9  => CPIX_NORMAL_INIT_58_BIT_09_C, 10 => CPIX_NORMAL_INIT_58_BIT_10_C, 11 => CPIX_NORMAL_INIT_58_BIT_11_C, 12 => CPIX_NORMAL_INIT_58_BIT_12_C, 13 => CPIX_NORMAL_INIT_58_BIT_13_C, 14 => CPIX_NORMAL_INIT_58_BIT_14_C);
   constant CPIX_NORMAL_INIT_59_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_59_BIT_00_C, 1  => CPIX_NORMAL_INIT_59_BIT_01_C, 2  => CPIX_NORMAL_INIT_59_BIT_02_C, 3  => CPIX_NORMAL_INIT_59_BIT_03_C, 4  => CPIX_NORMAL_INIT_59_BIT_04_C, 5  => CPIX_NORMAL_INIT_59_BIT_05_C, 6  => CPIX_NORMAL_INIT_59_BIT_06_C, 7  => CPIX_NORMAL_INIT_59_BIT_07_C, 8  => CPIX_NORMAL_INIT_59_BIT_08_C, 9  => CPIX_NORMAL_INIT_59_BIT_09_C, 10 => CPIX_NORMAL_INIT_59_BIT_10_C, 11 => CPIX_NORMAL_INIT_59_BIT_11_C, 12 => CPIX_NORMAL_INIT_59_BIT_12_C, 13 => CPIX_NORMAL_INIT_59_BIT_13_C, 14 => CPIX_NORMAL_INIT_59_BIT_14_C);
   constant CPIX_NORMAL_INIT_5A_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_5A_BIT_00_C, 1  => CPIX_NORMAL_INIT_5A_BIT_01_C, 2  => CPIX_NORMAL_INIT_5A_BIT_02_C, 3  => CPIX_NORMAL_INIT_5A_BIT_03_C, 4  => CPIX_NORMAL_INIT_5A_BIT_04_C, 5  => CPIX_NORMAL_INIT_5A_BIT_05_C, 6  => CPIX_NORMAL_INIT_5A_BIT_06_C, 7  => CPIX_NORMAL_INIT_5A_BIT_07_C, 8  => CPIX_NORMAL_INIT_5A_BIT_08_C, 9  => CPIX_NORMAL_INIT_5A_BIT_09_C, 10 => CPIX_NORMAL_INIT_5A_BIT_10_C, 11 => CPIX_NORMAL_INIT_5A_BIT_11_C, 12 => CPIX_NORMAL_INIT_5A_BIT_12_C, 13 => CPIX_NORMAL_INIT_5A_BIT_13_C, 14 => CPIX_NORMAL_INIT_5A_BIT_14_C);
   constant CPIX_NORMAL_INIT_5B_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_5B_BIT_00_C, 1  => CPIX_NORMAL_INIT_5B_BIT_01_C, 2  => CPIX_NORMAL_INIT_5B_BIT_02_C, 3  => CPIX_NORMAL_INIT_5B_BIT_03_C, 4  => CPIX_NORMAL_INIT_5B_BIT_04_C, 5  => CPIX_NORMAL_INIT_5B_BIT_05_C, 6  => CPIX_NORMAL_INIT_5B_BIT_06_C, 7  => CPIX_NORMAL_INIT_5B_BIT_07_C, 8  => CPIX_NORMAL_INIT_5B_BIT_08_C, 9  => CPIX_NORMAL_INIT_5B_BIT_09_C, 10 => CPIX_NORMAL_INIT_5B_BIT_10_C, 11 => CPIX_NORMAL_INIT_5B_BIT_11_C, 12 => CPIX_NORMAL_INIT_5B_BIT_12_C, 13 => CPIX_NORMAL_INIT_5B_BIT_13_C, 14 => CPIX_NORMAL_INIT_5B_BIT_14_C);
   constant CPIX_NORMAL_INIT_5C_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_5C_BIT_00_C, 1  => CPIX_NORMAL_INIT_5C_BIT_01_C, 2  => CPIX_NORMAL_INIT_5C_BIT_02_C, 3  => CPIX_NORMAL_INIT_5C_BIT_03_C, 4  => CPIX_NORMAL_INIT_5C_BIT_04_C, 5  => CPIX_NORMAL_INIT_5C_BIT_05_C, 6  => CPIX_NORMAL_INIT_5C_BIT_06_C, 7  => CPIX_NORMAL_INIT_5C_BIT_07_C, 8  => CPIX_NORMAL_INIT_5C_BIT_08_C, 9  => CPIX_NORMAL_INIT_5C_BIT_09_C, 10 => CPIX_NORMAL_INIT_5C_BIT_10_C, 11 => CPIX_NORMAL_INIT_5C_BIT_11_C, 12 => CPIX_NORMAL_INIT_5C_BIT_12_C, 13 => CPIX_NORMAL_INIT_5C_BIT_13_C, 14 => CPIX_NORMAL_INIT_5C_BIT_14_C);
   constant CPIX_NORMAL_INIT_5D_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_5D_BIT_00_C, 1  => CPIX_NORMAL_INIT_5D_BIT_01_C, 2  => CPIX_NORMAL_INIT_5D_BIT_02_C, 3  => CPIX_NORMAL_INIT_5D_BIT_03_C, 4  => CPIX_NORMAL_INIT_5D_BIT_04_C, 5  => CPIX_NORMAL_INIT_5D_BIT_05_C, 6  => CPIX_NORMAL_INIT_5D_BIT_06_C, 7  => CPIX_NORMAL_INIT_5D_BIT_07_C, 8  => CPIX_NORMAL_INIT_5D_BIT_08_C, 9  => CPIX_NORMAL_INIT_5D_BIT_09_C, 10 => CPIX_NORMAL_INIT_5D_BIT_10_C, 11 => CPIX_NORMAL_INIT_5D_BIT_11_C, 12 => CPIX_NORMAL_INIT_5D_BIT_12_C, 13 => CPIX_NORMAL_INIT_5D_BIT_13_C, 14 => CPIX_NORMAL_INIT_5D_BIT_14_C);
   constant CPIX_NORMAL_INIT_5E_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_5E_BIT_00_C, 1  => CPIX_NORMAL_INIT_5E_BIT_01_C, 2  => CPIX_NORMAL_INIT_5E_BIT_02_C, 3  => CPIX_NORMAL_INIT_5E_BIT_03_C, 4  => CPIX_NORMAL_INIT_5E_BIT_04_C, 5  => CPIX_NORMAL_INIT_5E_BIT_05_C, 6  => CPIX_NORMAL_INIT_5E_BIT_06_C, 7  => CPIX_NORMAL_INIT_5E_BIT_07_C, 8  => CPIX_NORMAL_INIT_5E_BIT_08_C, 9  => CPIX_NORMAL_INIT_5E_BIT_09_C, 10 => CPIX_NORMAL_INIT_5E_BIT_10_C, 11 => CPIX_NORMAL_INIT_5E_BIT_11_C, 12 => CPIX_NORMAL_INIT_5E_BIT_12_C, 13 => CPIX_NORMAL_INIT_5E_BIT_13_C, 14 => CPIX_NORMAL_INIT_5E_BIT_14_C);
   constant CPIX_NORMAL_INIT_5F_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_5F_BIT_00_C, 1  => CPIX_NORMAL_INIT_5F_BIT_01_C, 2  => CPIX_NORMAL_INIT_5F_BIT_02_C, 3  => CPIX_NORMAL_INIT_5F_BIT_03_C, 4  => CPIX_NORMAL_INIT_5F_BIT_04_C, 5  => CPIX_NORMAL_INIT_5F_BIT_05_C, 6  => CPIX_NORMAL_INIT_5F_BIT_06_C, 7  => CPIX_NORMAL_INIT_5F_BIT_07_C, 8  => CPIX_NORMAL_INIT_5F_BIT_08_C, 9  => CPIX_NORMAL_INIT_5F_BIT_09_C, 10 => CPIX_NORMAL_INIT_5F_BIT_10_C, 11 => CPIX_NORMAL_INIT_5F_BIT_11_C, 12 => CPIX_NORMAL_INIT_5F_BIT_12_C, 13 => CPIX_NORMAL_INIT_5F_BIT_13_C, 14 => CPIX_NORMAL_INIT_5F_BIT_14_C);
   constant CPIX_NORMAL_INIT_60_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_60_BIT_00_C, 1  => CPIX_NORMAL_INIT_60_BIT_01_C, 2  => CPIX_NORMAL_INIT_60_BIT_02_C, 3  => CPIX_NORMAL_INIT_60_BIT_03_C, 4  => CPIX_NORMAL_INIT_60_BIT_04_C, 5  => CPIX_NORMAL_INIT_60_BIT_05_C, 6  => CPIX_NORMAL_INIT_60_BIT_06_C, 7  => CPIX_NORMAL_INIT_60_BIT_07_C, 8  => CPIX_NORMAL_INIT_60_BIT_08_C, 9  => CPIX_NORMAL_INIT_60_BIT_09_C, 10 => CPIX_NORMAL_INIT_60_BIT_10_C, 11 => CPIX_NORMAL_INIT_60_BIT_11_C, 12 => CPIX_NORMAL_INIT_60_BIT_12_C, 13 => CPIX_NORMAL_INIT_60_BIT_13_C, 14 => CPIX_NORMAL_INIT_60_BIT_14_C);
   constant CPIX_NORMAL_INIT_61_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_61_BIT_00_C, 1  => CPIX_NORMAL_INIT_61_BIT_01_C, 2  => CPIX_NORMAL_INIT_61_BIT_02_C, 3  => CPIX_NORMAL_INIT_61_BIT_03_C, 4  => CPIX_NORMAL_INIT_61_BIT_04_C, 5  => CPIX_NORMAL_INIT_61_BIT_05_C, 6  => CPIX_NORMAL_INIT_61_BIT_06_C, 7  => CPIX_NORMAL_INIT_61_BIT_07_C, 8  => CPIX_NORMAL_INIT_61_BIT_08_C, 9  => CPIX_NORMAL_INIT_61_BIT_09_C, 10 => CPIX_NORMAL_INIT_61_BIT_10_C, 11 => CPIX_NORMAL_INIT_61_BIT_11_C, 12 => CPIX_NORMAL_INIT_61_BIT_12_C, 13 => CPIX_NORMAL_INIT_61_BIT_13_C, 14 => CPIX_NORMAL_INIT_61_BIT_14_C);
   constant CPIX_NORMAL_INIT_62_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_62_BIT_00_C, 1  => CPIX_NORMAL_INIT_62_BIT_01_C, 2  => CPIX_NORMAL_INIT_62_BIT_02_C, 3  => CPIX_NORMAL_INIT_62_BIT_03_C, 4  => CPIX_NORMAL_INIT_62_BIT_04_C, 5  => CPIX_NORMAL_INIT_62_BIT_05_C, 6  => CPIX_NORMAL_INIT_62_BIT_06_C, 7  => CPIX_NORMAL_INIT_62_BIT_07_C, 8  => CPIX_NORMAL_INIT_62_BIT_08_C, 9  => CPIX_NORMAL_INIT_62_BIT_09_C, 10 => CPIX_NORMAL_INIT_62_BIT_10_C, 11 => CPIX_NORMAL_INIT_62_BIT_11_C, 12 => CPIX_NORMAL_INIT_62_BIT_12_C, 13 => CPIX_NORMAL_INIT_62_BIT_13_C, 14 => CPIX_NORMAL_INIT_62_BIT_14_C);
   constant CPIX_NORMAL_INIT_63_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_63_BIT_00_C, 1  => CPIX_NORMAL_INIT_63_BIT_01_C, 2  => CPIX_NORMAL_INIT_63_BIT_02_C, 3  => CPIX_NORMAL_INIT_63_BIT_03_C, 4  => CPIX_NORMAL_INIT_63_BIT_04_C, 5  => CPIX_NORMAL_INIT_63_BIT_05_C, 6  => CPIX_NORMAL_INIT_63_BIT_06_C, 7  => CPIX_NORMAL_INIT_63_BIT_07_C, 8  => CPIX_NORMAL_INIT_63_BIT_08_C, 9  => CPIX_NORMAL_INIT_63_BIT_09_C, 10 => CPIX_NORMAL_INIT_63_BIT_10_C, 11 => CPIX_NORMAL_INIT_63_BIT_11_C, 12 => CPIX_NORMAL_INIT_63_BIT_12_C, 13 => CPIX_NORMAL_INIT_63_BIT_13_C, 14 => CPIX_NORMAL_INIT_63_BIT_14_C);
   constant CPIX_NORMAL_INIT_64_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_64_BIT_00_C, 1  => CPIX_NORMAL_INIT_64_BIT_01_C, 2  => CPIX_NORMAL_INIT_64_BIT_02_C, 3  => CPIX_NORMAL_INIT_64_BIT_03_C, 4  => CPIX_NORMAL_INIT_64_BIT_04_C, 5  => CPIX_NORMAL_INIT_64_BIT_05_C, 6  => CPIX_NORMAL_INIT_64_BIT_06_C, 7  => CPIX_NORMAL_INIT_64_BIT_07_C, 8  => CPIX_NORMAL_INIT_64_BIT_08_C, 9  => CPIX_NORMAL_INIT_64_BIT_09_C, 10 => CPIX_NORMAL_INIT_64_BIT_10_C, 11 => CPIX_NORMAL_INIT_64_BIT_11_C, 12 => CPIX_NORMAL_INIT_64_BIT_12_C, 13 => CPIX_NORMAL_INIT_64_BIT_13_C, 14 => CPIX_NORMAL_INIT_64_BIT_14_C);
   constant CPIX_NORMAL_INIT_65_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_65_BIT_00_C, 1  => CPIX_NORMAL_INIT_65_BIT_01_C, 2  => CPIX_NORMAL_INIT_65_BIT_02_C, 3  => CPIX_NORMAL_INIT_65_BIT_03_C, 4  => CPIX_NORMAL_INIT_65_BIT_04_C, 5  => CPIX_NORMAL_INIT_65_BIT_05_C, 6  => CPIX_NORMAL_INIT_65_BIT_06_C, 7  => CPIX_NORMAL_INIT_65_BIT_07_C, 8  => CPIX_NORMAL_INIT_65_BIT_08_C, 9  => CPIX_NORMAL_INIT_65_BIT_09_C, 10 => CPIX_NORMAL_INIT_65_BIT_10_C, 11 => CPIX_NORMAL_INIT_65_BIT_11_C, 12 => CPIX_NORMAL_INIT_65_BIT_12_C, 13 => CPIX_NORMAL_INIT_65_BIT_13_C, 14 => CPIX_NORMAL_INIT_65_BIT_14_C);
   constant CPIX_NORMAL_INIT_66_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_66_BIT_00_C, 1  => CPIX_NORMAL_INIT_66_BIT_01_C, 2  => CPIX_NORMAL_INIT_66_BIT_02_C, 3  => CPIX_NORMAL_INIT_66_BIT_03_C, 4  => CPIX_NORMAL_INIT_66_BIT_04_C, 5  => CPIX_NORMAL_INIT_66_BIT_05_C, 6  => CPIX_NORMAL_INIT_66_BIT_06_C, 7  => CPIX_NORMAL_INIT_66_BIT_07_C, 8  => CPIX_NORMAL_INIT_66_BIT_08_C, 9  => CPIX_NORMAL_INIT_66_BIT_09_C, 10 => CPIX_NORMAL_INIT_66_BIT_10_C, 11 => CPIX_NORMAL_INIT_66_BIT_11_C, 12 => CPIX_NORMAL_INIT_66_BIT_12_C, 13 => CPIX_NORMAL_INIT_66_BIT_13_C, 14 => CPIX_NORMAL_INIT_66_BIT_14_C);
   constant CPIX_NORMAL_INIT_67_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_67_BIT_00_C, 1  => CPIX_NORMAL_INIT_67_BIT_01_C, 2  => CPIX_NORMAL_INIT_67_BIT_02_C, 3  => CPIX_NORMAL_INIT_67_BIT_03_C, 4  => CPIX_NORMAL_INIT_67_BIT_04_C, 5  => CPIX_NORMAL_INIT_67_BIT_05_C, 6  => CPIX_NORMAL_INIT_67_BIT_06_C, 7  => CPIX_NORMAL_INIT_67_BIT_07_C, 8  => CPIX_NORMAL_INIT_67_BIT_08_C, 9  => CPIX_NORMAL_INIT_67_BIT_09_C, 10 => CPIX_NORMAL_INIT_67_BIT_10_C, 11 => CPIX_NORMAL_INIT_67_BIT_11_C, 12 => CPIX_NORMAL_INIT_67_BIT_12_C, 13 => CPIX_NORMAL_INIT_67_BIT_13_C, 14 => CPIX_NORMAL_INIT_67_BIT_14_C);
   constant CPIX_NORMAL_INIT_68_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_68_BIT_00_C, 1  => CPIX_NORMAL_INIT_68_BIT_01_C, 2  => CPIX_NORMAL_INIT_68_BIT_02_C, 3  => CPIX_NORMAL_INIT_68_BIT_03_C, 4  => CPIX_NORMAL_INIT_68_BIT_04_C, 5  => CPIX_NORMAL_INIT_68_BIT_05_C, 6  => CPIX_NORMAL_INIT_68_BIT_06_C, 7  => CPIX_NORMAL_INIT_68_BIT_07_C, 8  => CPIX_NORMAL_INIT_68_BIT_08_C, 9  => CPIX_NORMAL_INIT_68_BIT_09_C, 10 => CPIX_NORMAL_INIT_68_BIT_10_C, 11 => CPIX_NORMAL_INIT_68_BIT_11_C, 12 => CPIX_NORMAL_INIT_68_BIT_12_C, 13 => CPIX_NORMAL_INIT_68_BIT_13_C, 14 => CPIX_NORMAL_INIT_68_BIT_14_C);
   constant CPIX_NORMAL_INIT_69_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_69_BIT_00_C, 1  => CPIX_NORMAL_INIT_69_BIT_01_C, 2  => CPIX_NORMAL_INIT_69_BIT_02_C, 3  => CPIX_NORMAL_INIT_69_BIT_03_C, 4  => CPIX_NORMAL_INIT_69_BIT_04_C, 5  => CPIX_NORMAL_INIT_69_BIT_05_C, 6  => CPIX_NORMAL_INIT_69_BIT_06_C, 7  => CPIX_NORMAL_INIT_69_BIT_07_C, 8  => CPIX_NORMAL_INIT_69_BIT_08_C, 9  => CPIX_NORMAL_INIT_69_BIT_09_C, 10 => CPIX_NORMAL_INIT_69_BIT_10_C, 11 => CPIX_NORMAL_INIT_69_BIT_11_C, 12 => CPIX_NORMAL_INIT_69_BIT_12_C, 13 => CPIX_NORMAL_INIT_69_BIT_13_C, 14 => CPIX_NORMAL_INIT_69_BIT_14_C);
   constant CPIX_NORMAL_INIT_6A_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_6A_BIT_00_C, 1  => CPIX_NORMAL_INIT_6A_BIT_01_C, 2  => CPIX_NORMAL_INIT_6A_BIT_02_C, 3  => CPIX_NORMAL_INIT_6A_BIT_03_C, 4  => CPIX_NORMAL_INIT_6A_BIT_04_C, 5  => CPIX_NORMAL_INIT_6A_BIT_05_C, 6  => CPIX_NORMAL_INIT_6A_BIT_06_C, 7  => CPIX_NORMAL_INIT_6A_BIT_07_C, 8  => CPIX_NORMAL_INIT_6A_BIT_08_C, 9  => CPIX_NORMAL_INIT_6A_BIT_09_C, 10 => CPIX_NORMAL_INIT_6A_BIT_10_C, 11 => CPIX_NORMAL_INIT_6A_BIT_11_C, 12 => CPIX_NORMAL_INIT_6A_BIT_12_C, 13 => CPIX_NORMAL_INIT_6A_BIT_13_C, 14 => CPIX_NORMAL_INIT_6A_BIT_14_C);
   constant CPIX_NORMAL_INIT_6B_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_6B_BIT_00_C, 1  => CPIX_NORMAL_INIT_6B_BIT_01_C, 2  => CPIX_NORMAL_INIT_6B_BIT_02_C, 3  => CPIX_NORMAL_INIT_6B_BIT_03_C, 4  => CPIX_NORMAL_INIT_6B_BIT_04_C, 5  => CPIX_NORMAL_INIT_6B_BIT_05_C, 6  => CPIX_NORMAL_INIT_6B_BIT_06_C, 7  => CPIX_NORMAL_INIT_6B_BIT_07_C, 8  => CPIX_NORMAL_INIT_6B_BIT_08_C, 9  => CPIX_NORMAL_INIT_6B_BIT_09_C, 10 => CPIX_NORMAL_INIT_6B_BIT_10_C, 11 => CPIX_NORMAL_INIT_6B_BIT_11_C, 12 => CPIX_NORMAL_INIT_6B_BIT_12_C, 13 => CPIX_NORMAL_INIT_6B_BIT_13_C, 14 => CPIX_NORMAL_INIT_6B_BIT_14_C);
   constant CPIX_NORMAL_INIT_6C_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_6C_BIT_00_C, 1  => CPIX_NORMAL_INIT_6C_BIT_01_C, 2  => CPIX_NORMAL_INIT_6C_BIT_02_C, 3  => CPIX_NORMAL_INIT_6C_BIT_03_C, 4  => CPIX_NORMAL_INIT_6C_BIT_04_C, 5  => CPIX_NORMAL_INIT_6C_BIT_05_C, 6  => CPIX_NORMAL_INIT_6C_BIT_06_C, 7  => CPIX_NORMAL_INIT_6C_BIT_07_C, 8  => CPIX_NORMAL_INIT_6C_BIT_08_C, 9  => CPIX_NORMAL_INIT_6C_BIT_09_C, 10 => CPIX_NORMAL_INIT_6C_BIT_10_C, 11 => CPIX_NORMAL_INIT_6C_BIT_11_C, 12 => CPIX_NORMAL_INIT_6C_BIT_12_C, 13 => CPIX_NORMAL_INIT_6C_BIT_13_C, 14 => CPIX_NORMAL_INIT_6C_BIT_14_C);
   constant CPIX_NORMAL_INIT_6D_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_6D_BIT_00_C, 1  => CPIX_NORMAL_INIT_6D_BIT_01_C, 2  => CPIX_NORMAL_INIT_6D_BIT_02_C, 3  => CPIX_NORMAL_INIT_6D_BIT_03_C, 4  => CPIX_NORMAL_INIT_6D_BIT_04_C, 5  => CPIX_NORMAL_INIT_6D_BIT_05_C, 6  => CPIX_NORMAL_INIT_6D_BIT_06_C, 7  => CPIX_NORMAL_INIT_6D_BIT_07_C, 8  => CPIX_NORMAL_INIT_6D_BIT_08_C, 9  => CPIX_NORMAL_INIT_6D_BIT_09_C, 10 => CPIX_NORMAL_INIT_6D_BIT_10_C, 11 => CPIX_NORMAL_INIT_6D_BIT_11_C, 12 => CPIX_NORMAL_INIT_6D_BIT_12_C, 13 => CPIX_NORMAL_INIT_6D_BIT_13_C, 14 => CPIX_NORMAL_INIT_6D_BIT_14_C);
   constant CPIX_NORMAL_INIT_6E_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_6E_BIT_00_C, 1  => CPIX_NORMAL_INIT_6E_BIT_01_C, 2  => CPIX_NORMAL_INIT_6E_BIT_02_C, 3  => CPIX_NORMAL_INIT_6E_BIT_03_C, 4  => CPIX_NORMAL_INIT_6E_BIT_04_C, 5  => CPIX_NORMAL_INIT_6E_BIT_05_C, 6  => CPIX_NORMAL_INIT_6E_BIT_06_C, 7  => CPIX_NORMAL_INIT_6E_BIT_07_C, 8  => CPIX_NORMAL_INIT_6E_BIT_08_C, 9  => CPIX_NORMAL_INIT_6E_BIT_09_C, 10 => CPIX_NORMAL_INIT_6E_BIT_10_C, 11 => CPIX_NORMAL_INIT_6E_BIT_11_C, 12 => CPIX_NORMAL_INIT_6E_BIT_12_C, 13 => CPIX_NORMAL_INIT_6E_BIT_13_C, 14 => CPIX_NORMAL_INIT_6E_BIT_14_C);
   constant CPIX_NORMAL_INIT_6F_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_6F_BIT_00_C, 1  => CPIX_NORMAL_INIT_6F_BIT_01_C, 2  => CPIX_NORMAL_INIT_6F_BIT_02_C, 3  => CPIX_NORMAL_INIT_6F_BIT_03_C, 4  => CPIX_NORMAL_INIT_6F_BIT_04_C, 5  => CPIX_NORMAL_INIT_6F_BIT_05_C, 6  => CPIX_NORMAL_INIT_6F_BIT_06_C, 7  => CPIX_NORMAL_INIT_6F_BIT_07_C, 8  => CPIX_NORMAL_INIT_6F_BIT_08_C, 9  => CPIX_NORMAL_INIT_6F_BIT_09_C, 10 => CPIX_NORMAL_INIT_6F_BIT_10_C, 11 => CPIX_NORMAL_INIT_6F_BIT_11_C, 12 => CPIX_NORMAL_INIT_6F_BIT_12_C, 13 => CPIX_NORMAL_INIT_6F_BIT_13_C, 14 => CPIX_NORMAL_INIT_6F_BIT_14_C);
   constant CPIX_NORMAL_INIT_70_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_70_BIT_00_C, 1  => CPIX_NORMAL_INIT_70_BIT_01_C, 2  => CPIX_NORMAL_INIT_70_BIT_02_C, 3  => CPIX_NORMAL_INIT_70_BIT_03_C, 4  => CPIX_NORMAL_INIT_70_BIT_04_C, 5  => CPIX_NORMAL_INIT_70_BIT_05_C, 6  => CPIX_NORMAL_INIT_70_BIT_06_C, 7  => CPIX_NORMAL_INIT_70_BIT_07_C, 8  => CPIX_NORMAL_INIT_70_BIT_08_C, 9  => CPIX_NORMAL_INIT_70_BIT_09_C, 10 => CPIX_NORMAL_INIT_70_BIT_10_C, 11 => CPIX_NORMAL_INIT_70_BIT_11_C, 12 => CPIX_NORMAL_INIT_70_BIT_12_C, 13 => CPIX_NORMAL_INIT_70_BIT_13_C, 14 => CPIX_NORMAL_INIT_70_BIT_14_C);
   constant CPIX_NORMAL_INIT_71_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_71_BIT_00_C, 1  => CPIX_NORMAL_INIT_71_BIT_01_C, 2  => CPIX_NORMAL_INIT_71_BIT_02_C, 3  => CPIX_NORMAL_INIT_71_BIT_03_C, 4  => CPIX_NORMAL_INIT_71_BIT_04_C, 5  => CPIX_NORMAL_INIT_71_BIT_05_C, 6  => CPIX_NORMAL_INIT_71_BIT_06_C, 7  => CPIX_NORMAL_INIT_71_BIT_07_C, 8  => CPIX_NORMAL_INIT_71_BIT_08_C, 9  => CPIX_NORMAL_INIT_71_BIT_09_C, 10 => CPIX_NORMAL_INIT_71_BIT_10_C, 11 => CPIX_NORMAL_INIT_71_BIT_11_C, 12 => CPIX_NORMAL_INIT_71_BIT_12_C, 13 => CPIX_NORMAL_INIT_71_BIT_13_C, 14 => CPIX_NORMAL_INIT_71_BIT_14_C);
   constant CPIX_NORMAL_INIT_72_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_72_BIT_00_C, 1  => CPIX_NORMAL_INIT_72_BIT_01_C, 2  => CPIX_NORMAL_INIT_72_BIT_02_C, 3  => CPIX_NORMAL_INIT_72_BIT_03_C, 4  => CPIX_NORMAL_INIT_72_BIT_04_C, 5  => CPIX_NORMAL_INIT_72_BIT_05_C, 6  => CPIX_NORMAL_INIT_72_BIT_06_C, 7  => CPIX_NORMAL_INIT_72_BIT_07_C, 8  => CPIX_NORMAL_INIT_72_BIT_08_C, 9  => CPIX_NORMAL_INIT_72_BIT_09_C, 10 => CPIX_NORMAL_INIT_72_BIT_10_C, 11 => CPIX_NORMAL_INIT_72_BIT_11_C, 12 => CPIX_NORMAL_INIT_72_BIT_12_C, 13 => CPIX_NORMAL_INIT_72_BIT_13_C, 14 => CPIX_NORMAL_INIT_72_BIT_14_C);
   constant CPIX_NORMAL_INIT_73_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_73_BIT_00_C, 1  => CPIX_NORMAL_INIT_73_BIT_01_C, 2  => CPIX_NORMAL_INIT_73_BIT_02_C, 3  => CPIX_NORMAL_INIT_73_BIT_03_C, 4  => CPIX_NORMAL_INIT_73_BIT_04_C, 5  => CPIX_NORMAL_INIT_73_BIT_05_C, 6  => CPIX_NORMAL_INIT_73_BIT_06_C, 7  => CPIX_NORMAL_INIT_73_BIT_07_C, 8  => CPIX_NORMAL_INIT_73_BIT_08_C, 9  => CPIX_NORMAL_INIT_73_BIT_09_C, 10 => CPIX_NORMAL_INIT_73_BIT_10_C, 11 => CPIX_NORMAL_INIT_73_BIT_11_C, 12 => CPIX_NORMAL_INIT_73_BIT_12_C, 13 => CPIX_NORMAL_INIT_73_BIT_13_C, 14 => CPIX_NORMAL_INIT_73_BIT_14_C);
   constant CPIX_NORMAL_INIT_74_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_74_BIT_00_C, 1  => CPIX_NORMAL_INIT_74_BIT_01_C, 2  => CPIX_NORMAL_INIT_74_BIT_02_C, 3  => CPIX_NORMAL_INIT_74_BIT_03_C, 4  => CPIX_NORMAL_INIT_74_BIT_04_C, 5  => CPIX_NORMAL_INIT_74_BIT_05_C, 6  => CPIX_NORMAL_INIT_74_BIT_06_C, 7  => CPIX_NORMAL_INIT_74_BIT_07_C, 8  => CPIX_NORMAL_INIT_74_BIT_08_C, 9  => CPIX_NORMAL_INIT_74_BIT_09_C, 10 => CPIX_NORMAL_INIT_74_BIT_10_C, 11 => CPIX_NORMAL_INIT_74_BIT_11_C, 12 => CPIX_NORMAL_INIT_74_BIT_12_C, 13 => CPIX_NORMAL_INIT_74_BIT_13_C, 14 => CPIX_NORMAL_INIT_74_BIT_14_C);
   constant CPIX_NORMAL_INIT_75_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_75_BIT_00_C, 1  => CPIX_NORMAL_INIT_75_BIT_01_C, 2  => CPIX_NORMAL_INIT_75_BIT_02_C, 3  => CPIX_NORMAL_INIT_75_BIT_03_C, 4  => CPIX_NORMAL_INIT_75_BIT_04_C, 5  => CPIX_NORMAL_INIT_75_BIT_05_C, 6  => CPIX_NORMAL_INIT_75_BIT_06_C, 7  => CPIX_NORMAL_INIT_75_BIT_07_C, 8  => CPIX_NORMAL_INIT_75_BIT_08_C, 9  => CPIX_NORMAL_INIT_75_BIT_09_C, 10 => CPIX_NORMAL_INIT_75_BIT_10_C, 11 => CPIX_NORMAL_INIT_75_BIT_11_C, 12 => CPIX_NORMAL_INIT_75_BIT_12_C, 13 => CPIX_NORMAL_INIT_75_BIT_13_C, 14 => CPIX_NORMAL_INIT_75_BIT_14_C);
   constant CPIX_NORMAL_INIT_76_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_76_BIT_00_C, 1  => CPIX_NORMAL_INIT_76_BIT_01_C, 2  => CPIX_NORMAL_INIT_76_BIT_02_C, 3  => CPIX_NORMAL_INIT_76_BIT_03_C, 4  => CPIX_NORMAL_INIT_76_BIT_04_C, 5  => CPIX_NORMAL_INIT_76_BIT_05_C, 6  => CPIX_NORMAL_INIT_76_BIT_06_C, 7  => CPIX_NORMAL_INIT_76_BIT_07_C, 8  => CPIX_NORMAL_INIT_76_BIT_08_C, 9  => CPIX_NORMAL_INIT_76_BIT_09_C, 10 => CPIX_NORMAL_INIT_76_BIT_10_C, 11 => CPIX_NORMAL_INIT_76_BIT_11_C, 12 => CPIX_NORMAL_INIT_76_BIT_12_C, 13 => CPIX_NORMAL_INIT_76_BIT_13_C, 14 => CPIX_NORMAL_INIT_76_BIT_14_C);
   constant CPIX_NORMAL_INIT_77_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_77_BIT_00_C, 1  => CPIX_NORMAL_INIT_77_BIT_01_C, 2  => CPIX_NORMAL_INIT_77_BIT_02_C, 3  => CPIX_NORMAL_INIT_77_BIT_03_C, 4  => CPIX_NORMAL_INIT_77_BIT_04_C, 5  => CPIX_NORMAL_INIT_77_BIT_05_C, 6  => CPIX_NORMAL_INIT_77_BIT_06_C, 7  => CPIX_NORMAL_INIT_77_BIT_07_C, 8  => CPIX_NORMAL_INIT_77_BIT_08_C, 9  => CPIX_NORMAL_INIT_77_BIT_09_C, 10 => CPIX_NORMAL_INIT_77_BIT_10_C, 11 => CPIX_NORMAL_INIT_77_BIT_11_C, 12 => CPIX_NORMAL_INIT_77_BIT_12_C, 13 => CPIX_NORMAL_INIT_77_BIT_13_C, 14 => CPIX_NORMAL_INIT_77_BIT_14_C);
   constant CPIX_NORMAL_INIT_78_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_78_BIT_00_C, 1  => CPIX_NORMAL_INIT_78_BIT_01_C, 2  => CPIX_NORMAL_INIT_78_BIT_02_C, 3  => CPIX_NORMAL_INIT_78_BIT_03_C, 4  => CPIX_NORMAL_INIT_78_BIT_04_C, 5  => CPIX_NORMAL_INIT_78_BIT_05_C, 6  => CPIX_NORMAL_INIT_78_BIT_06_C, 7  => CPIX_NORMAL_INIT_78_BIT_07_C, 8  => CPIX_NORMAL_INIT_78_BIT_08_C, 9  => CPIX_NORMAL_INIT_78_BIT_09_C, 10 => CPIX_NORMAL_INIT_78_BIT_10_C, 11 => CPIX_NORMAL_INIT_78_BIT_11_C, 12 => CPIX_NORMAL_INIT_78_BIT_12_C, 13 => CPIX_NORMAL_INIT_78_BIT_13_C, 14 => CPIX_NORMAL_INIT_78_BIT_14_C);
   constant CPIX_NORMAL_INIT_79_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_79_BIT_00_C, 1  => CPIX_NORMAL_INIT_79_BIT_01_C, 2  => CPIX_NORMAL_INIT_79_BIT_02_C, 3  => CPIX_NORMAL_INIT_79_BIT_03_C, 4  => CPIX_NORMAL_INIT_79_BIT_04_C, 5  => CPIX_NORMAL_INIT_79_BIT_05_C, 6  => CPIX_NORMAL_INIT_79_BIT_06_C, 7  => CPIX_NORMAL_INIT_79_BIT_07_C, 8  => CPIX_NORMAL_INIT_79_BIT_08_C, 9  => CPIX_NORMAL_INIT_79_BIT_09_C, 10 => CPIX_NORMAL_INIT_79_BIT_10_C, 11 => CPIX_NORMAL_INIT_79_BIT_11_C, 12 => CPIX_NORMAL_INIT_79_BIT_12_C, 13 => CPIX_NORMAL_INIT_79_BIT_13_C, 14 => CPIX_NORMAL_INIT_79_BIT_14_C);
   constant CPIX_NORMAL_INIT_7A_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_7A_BIT_00_C, 1  => CPIX_NORMAL_INIT_7A_BIT_01_C, 2  => CPIX_NORMAL_INIT_7A_BIT_02_C, 3  => CPIX_NORMAL_INIT_7A_BIT_03_C, 4  => CPIX_NORMAL_INIT_7A_BIT_04_C, 5  => CPIX_NORMAL_INIT_7A_BIT_05_C, 6  => CPIX_NORMAL_INIT_7A_BIT_06_C, 7  => CPIX_NORMAL_INIT_7A_BIT_07_C, 8  => CPIX_NORMAL_INIT_7A_BIT_08_C, 9  => CPIX_NORMAL_INIT_7A_BIT_09_C, 10 => CPIX_NORMAL_INIT_7A_BIT_10_C, 11 => CPIX_NORMAL_INIT_7A_BIT_11_C, 12 => CPIX_NORMAL_INIT_7A_BIT_12_C, 13 => CPIX_NORMAL_INIT_7A_BIT_13_C, 14 => CPIX_NORMAL_INIT_7A_BIT_14_C);
   constant CPIX_NORMAL_INIT_7B_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_7B_BIT_00_C, 1  => CPIX_NORMAL_INIT_7B_BIT_01_C, 2  => CPIX_NORMAL_INIT_7B_BIT_02_C, 3  => CPIX_NORMAL_INIT_7B_BIT_03_C, 4  => CPIX_NORMAL_INIT_7B_BIT_04_C, 5  => CPIX_NORMAL_INIT_7B_BIT_05_C, 6  => CPIX_NORMAL_INIT_7B_BIT_06_C, 7  => CPIX_NORMAL_INIT_7B_BIT_07_C, 8  => CPIX_NORMAL_INIT_7B_BIT_08_C, 9  => CPIX_NORMAL_INIT_7B_BIT_09_C, 10 => CPIX_NORMAL_INIT_7B_BIT_10_C, 11 => CPIX_NORMAL_INIT_7B_BIT_11_C, 12 => CPIX_NORMAL_INIT_7B_BIT_12_C, 13 => CPIX_NORMAL_INIT_7B_BIT_13_C, 14 => CPIX_NORMAL_INIT_7B_BIT_14_C);
   constant CPIX_NORMAL_INIT_7C_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_7C_BIT_00_C, 1  => CPIX_NORMAL_INIT_7C_BIT_01_C, 2  => CPIX_NORMAL_INIT_7C_BIT_02_C, 3  => CPIX_NORMAL_INIT_7C_BIT_03_C, 4  => CPIX_NORMAL_INIT_7C_BIT_04_C, 5  => CPIX_NORMAL_INIT_7C_BIT_05_C, 6  => CPIX_NORMAL_INIT_7C_BIT_06_C, 7  => CPIX_NORMAL_INIT_7C_BIT_07_C, 8  => CPIX_NORMAL_INIT_7C_BIT_08_C, 9  => CPIX_NORMAL_INIT_7C_BIT_09_C, 10 => CPIX_NORMAL_INIT_7C_BIT_10_C, 11 => CPIX_NORMAL_INIT_7C_BIT_11_C, 12 => CPIX_NORMAL_INIT_7C_BIT_12_C, 13 => CPIX_NORMAL_INIT_7C_BIT_13_C, 14 => CPIX_NORMAL_INIT_7C_BIT_14_C);
   constant CPIX_NORMAL_INIT_7D_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_7D_BIT_00_C, 1  => CPIX_NORMAL_INIT_7D_BIT_01_C, 2  => CPIX_NORMAL_INIT_7D_BIT_02_C, 3  => CPIX_NORMAL_INIT_7D_BIT_03_C, 4  => CPIX_NORMAL_INIT_7D_BIT_04_C, 5  => CPIX_NORMAL_INIT_7D_BIT_05_C, 6  => CPIX_NORMAL_INIT_7D_BIT_06_C, 7  => CPIX_NORMAL_INIT_7D_BIT_07_C, 8  => CPIX_NORMAL_INIT_7D_BIT_08_C, 9  => CPIX_NORMAL_INIT_7D_BIT_09_C, 10 => CPIX_NORMAL_INIT_7D_BIT_10_C, 11 => CPIX_NORMAL_INIT_7D_BIT_11_C, 12 => CPIX_NORMAL_INIT_7D_BIT_12_C, 13 => CPIX_NORMAL_INIT_7D_BIT_13_C, 14 => CPIX_NORMAL_INIT_7D_BIT_14_C);
   constant CPIX_NORMAL_INIT_7E_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_7E_BIT_00_C, 1  => CPIX_NORMAL_INIT_7E_BIT_01_C, 2  => CPIX_NORMAL_INIT_7E_BIT_02_C, 3  => CPIX_NORMAL_INIT_7E_BIT_03_C, 4  => CPIX_NORMAL_INIT_7E_BIT_04_C, 5  => CPIX_NORMAL_INIT_7E_BIT_05_C, 6  => CPIX_NORMAL_INIT_7E_BIT_06_C, 7  => CPIX_NORMAL_INIT_7E_BIT_07_C, 8  => CPIX_NORMAL_INIT_7E_BIT_08_C, 9  => CPIX_NORMAL_INIT_7E_BIT_09_C, 10 => CPIX_NORMAL_INIT_7E_BIT_10_C, 11 => CPIX_NORMAL_INIT_7E_BIT_11_C, 12 => CPIX_NORMAL_INIT_7E_BIT_12_C, 13 => CPIX_NORMAL_INIT_7E_BIT_13_C, 14 => CPIX_NORMAL_INIT_7E_BIT_14_C);
   constant CPIX_NORMAL_INIT_7F_BITS_C : Bit256Array(14 downto 0) := (0  => CPIX_NORMAL_INIT_7F_BIT_00_C, 1  => CPIX_NORMAL_INIT_7F_BIT_01_C, 2  => CPIX_NORMAL_INIT_7F_BIT_02_C, 3  => CPIX_NORMAL_INIT_7F_BIT_03_C, 4  => CPIX_NORMAL_INIT_7F_BIT_04_C, 5  => CPIX_NORMAL_INIT_7F_BIT_05_C, 6  => CPIX_NORMAL_INIT_7F_BIT_06_C, 7  => CPIX_NORMAL_INIT_7F_BIT_07_C, 8  => CPIX_NORMAL_INIT_7F_BIT_08_C, 9  => CPIX_NORMAL_INIT_7F_BIT_09_C, 10 => CPIX_NORMAL_INIT_7F_BIT_10_C, 11 => CPIX_NORMAL_INIT_7F_BIT_11_C, 12 => CPIX_NORMAL_INIT_7F_BIT_12_C, 13 => CPIX_NORMAL_INIT_7F_BIT_13_C, 14 => CPIX_NORMAL_INIT_7F_BIT_14_C);



end CpixLUTPkg;
