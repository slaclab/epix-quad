../code/EpixStartupCode.vhd